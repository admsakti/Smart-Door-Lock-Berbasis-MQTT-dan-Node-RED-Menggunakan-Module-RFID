PK   {c�Xx��\�  oa    cirkitFile.json�]Y�G��+������Z��k����A�:-�l�e����Qų�$�Ivc�z���2##3����*����_��y�\��_���by?y��t�%]_�㿲��aq?_/�?�҇/��Կ'���$[�i�-�ϼ(t�s�'�y��Lg�,����z�UZ�ٜM�~��?���C�|����_�K�}���i���NR_�$�Y�K��RUs=�<��}��a���*�OJ/8�u�xQ%��*l��&�s9̹�yU$ާ2Q����T&K�7o��d�I�憴plΉ�·�.K����B���˝N��9/R�:��/m�9i�a�m��Ʋ�WY�&��Q���FKL��,��T�%.��~�-;����@������G�J���*6�d��ܑy�R`sO�Jt#3A&\p:T�]Y�I��<!sAח��0�$���$�`��5ly(U�R�q[)eU���dI�)�ei�S�Bv�+�7�%<�`��N���ڂr��R>�`.^n�	��f��&i�,8y�iX�*K
�L��L��9�H�M��*S08>vFٚ]}8�T�u�j��ݻ�cd��̏��֑ݻ����]�bdwP(qc����(g�PF�!W%f�I�C�R˜44QȚ��)�+r�2���U���( m͉��wݍ��C*5u҆���@m8�$!��6kA��5A<���S\��1�-��2�i�!J� 6��O����$͡���O2X�e^1����T�H�GSF�wVri�K���b�xn��d�U4^)H���"ds!c��9��v*aގ22mڌ6mA<����
�]Q���l![�V�GF��li����-���v!i$S��44-?�)CӴCX##S���%���+�E�O��Ъ#C�W�8�ҤX!ci5Tzhɑ'��T��q�e�C1�J:�޸XE�Bv=���:��PC��_diM/�x9�� 2a�ߌu]?��/n˗w���m�k��Rh�5��䛪�s�PSg�"j
��p�PS6��H��"�8E"Ԕ��(���(G�5�Fq8�D�)>��Q$B�R�8,Ţ�)L��S$J�2�H<E��<��EiS���hڛGS߱(mʛ"��4�~&�������@%���5�p3��&���:��f�ө'Qٞc�Tu�rƌ��i��K�\I!�!�|A�ɐ�rA��i� -��<P)�.숱6��2���c��h�ũ��BP�l}��T��֪����X�Q�"�[E���ᄮ{�|�i�H�O�A����,a�M�t�Ї-1�y1������m6�z]�)���%6���6?��V��*t `SާQ�M_�6#�����MHG�rv����Ӈ66U|���f}OK 6}{z]�y�T�Z����i^�)��'6[yZ{c3��56�xڌ�&O�T���i��;m&b3n��M�E�b�y��l�^3[��t]FHlݗO�UzGOlE ����p��&���H�6��(E"�IlE�(�Mb+
G�m[Q8�Dh�؊�Q$B��V�"�$��p��6�GE�����v4�ͣ)�X����8<E��<��Ei�؊�S4�ͣ)��[t*y� �E����-:� n.Hlѩ��[t*�s��V2q�R�$�"�����$��L�8 �qP,�XD��qP,�X�A���b�"�E��(F'��T�b�آS9�:�E������Nlѩ�ltb�$tb�N���[t*g��آS9�.�����uA'��Tή:�E�r�tb�N�</���J^�b�آS9�wщ-:���:�����~�m�y_k�(~�����Ū|�?ܥyY����(W��	o�9j����_:�z�����Ĝe��G�/ɟW>���2�}G~י:���9�e_Zy�O2�=� #M)j��Z��\VZn�5,QN�e%���֢b�Z�С�J�д���Ђ6�&M<U0C�hCʍPCk�pQ�<�1N>�H9���/`_���V(N_��ɧٍOS}������� ���:%����##Ԕ��x�~����AJ��:����O���Z�O�S��J)< �vH���̱4т��b��aRpT�e�'Z����iC�nɃ�F�(�)ׁ��=ʷ�I�k���o��w��_-����Z�!F�<�C���"�C��I"�C�����CS� ��~� �#�L�|��7�pJh��D���8%�Gv�C��\��mb\�p����%E�*�2�g"��A589�@�w�*��%�_����M�NW�Qʛ)q���䔈���Uh�$Z� {%�5<]Z\Y�F*����I�o���]1ƪ�e�kY���b�0�#0	���?k�� �/ֈ���:J7&��|��Ib���kH�����,�� }���[	b]�5w[^����l�o�E���Xs�b�M�s�X�����b=N�e98 V�D���� ��Z���7�9*wN�ŭ
x"����
L\~^�/^�#װ�.��y�r5F�����[��d��G'�ER���FZ9]S�*R��qdu�ɤ�5�B��ܢ^+�T˶���VoE�p�E\8��r�d�%]�D#��봽p���z�"�:��o\iF\Rl����7xHWM�H8���]/
����^[H�A�\�" �d-�PjI������"�z�Pla��b���L:�2M:�&m� �nF�N�%�8x�����:���1lyg��jd�щf�U�A�w�j�yT��y�>�z/�ٽŃ�����V74��s[�6�Pư�p��b�L��ڈ�7����QNI��pE0�m�k��h�Hux:����]��{*�%���ά�-ޗ	� 2�Nzg�$
o��?� ���r�śKW�y��Q*ϗ��rߧ
/���-
�o_q�3F�d<_�o��������������]��%�O�"������[\���:Io���7�tΩo�Il��$rA&��������
N"d�k7�\�Il��$rA&��^�����JM"d�k4�l�il�Τ�A���.��G�#�P:��T>"hQA��il���k��%9�t�I�Xӏؿ���%Z��F; ���srt΄����*3@�{褔��]��:*=z��W*|�Q��y�I_��[0ꋒ4�T��q6�� �Ie��(�r�m$�6�>=�	�T.�:\�:P0�-x��Կa�B�`��E�o�쐣���#�)��4q���X�C��~X;��Q�P�L�	݀�v�3��nF߿��-�"���fF��X,�]���xS}g�Z@���rv�����'7�:qk���3"9�Ռ����6���ᄾֳ3� ���{v�����Z_�?;�ho�a�����}h@�����}h�Z�WF_�Y{_�z �(�����o�o��㤞b��j�ւP�@��v5��mT�[�Ӎ-� ���xl�Fa�=�;4�c�_�]�[S0���5�RM~�y����es��c����c��`��>��#����9b�j�Fӵ; {\�jJ	ۤ�"�U�\�)����,MY����#��˘w2)����%�pU薖�	^nZf��	�,1֤�7���%��JXǼ����4Rj�\�X$*S��'�;��H������8,�`0zf�$�+��)�Z�٦%`�`(J�<2^���$��`��ߴ4�����VR��d�2Ɍ��U������i�j�Y�2Q��o�JX��*`Nlifʋ�Þ�,y�~J+3��*�kx�����V�M���{��_Q"����x��G1�)�!�r#�:)~%����qK.�x��0%T@����h����+��s#I�Po�[n���涨�OY�R}���N���D�z�T��pC�y�6�pC���pC�$���$�z�H?�<��M. �G+s�;I��3�kJ���afnrsI?T=��m.���#���I���YZ����wiV��>SG������7��;O���?�G��Hn�ޣ&+���g;>� #j�L���#�d��L���>r�G;�,�ڱyd���V|�V��X|�X|`�v���i�ݴy�|7o�0���͏|��}���-�54���Z&������V
�/K���rn�\���z*�±�b�3��w.[��>@8c�E��2�Ӳ�K��*����?�gņ�;�@���#�Ruma�F:L�Fu/n�ߥ�:��G����C�Z/�&V���}��Z>a�׫���0��������t�kz�T���~�_ s�����������۪f >��������mU���bU��kXE��_���*��O��������\�{�V��������S�&B�
�zX>.֋%��G����@p+7���ڙ��	���	K\s�=��deU(��9��ZM&Z��S[�B[&m����T����t��\����*;�,a���t��d���˺&�X�w�v�?r��L���t���3���l�_]�\���XX?�垳	�ə��Mg���3��p[�S���ύ��˔�*���%i&A�W�J��)*����͈̠�	K�.S��z�_%�,��*m~Ѯs�,��������%�GR�zJ㥃^Vʹ�����4�^�J�v@j�`��SPBk�o ]� �c���3.$s~_?���83�ڪ�㝪
VȬЉ����� �%lW�:+gV���*M�ݩ��³�!�6pvf�%�ܑ.��P���0�h�Yf��r3��n{8��J�4=�W	H(=�,)S8Sxj��r�r��4*K�]��9�Z'[�R�H���Z��6Q[�2��ki�;v�x�K����.Z�Q�����DZ#^�1��j�0��g� ��4�na�T*9^�=����Da%/x�[]%��O�UIU���܈��<�/T2�/D��KpP�Lm~�>t����8n6���b���Й-%/e�k�&��U�;_�-�e���,N�r�\�.�hpq���6�ƽ l��D�l�j��=����fX�[�(OG���2S������%�É�E���<PP�j�mj�J6`����lg�\X�_`���kqت�|x/��M˻t�X�~Dw��=壿lI�9ݓ[�h:���v��~��c���~?v��Ϻ�"��ϫ��}�ny�<灙n��t����'|����4o�|h�]��0�$�:�������;�u��_X�����'*�YjAJG��[>�Wo���z����!6� ���y����j���g�L'�t�X��v,@���������I��*�{�U8S�q^��L8x�ݛ�Ż7���*��2zS�F̘_\
���ZM��W�)m���}�FRT��Kҿ|W�9�<]7�x��W)������N	˝�LN�c3a��I��������J_���z����z����W���j~�3�I	��T)?�`�x��˫H(���I臧�����p�ӛ�޽
髐�� �ZϤ�{f�1�O-�3�����(������)�IRZޕ��EQ�髐�
�m��ș3�Q���v���i��`J(Ϯ6B�W�D�����r���|��X�_^��UJo+�`�r�,�hB9e�T���
m�WҸ��)ꭶ$��]ޥ��J�t�T:Af�	p���vj�9pB�u �^����I_�p����^e�U6o)�N��3�����iµ�9Ƽs�K.��N����u�����3qT��	�F��P��e,箰��>K�ȫ�e�%E�<������t5Q@jz&�����_�JC�Զbөó�>�1�-�����6�8�aW����^���:��g���>��n���PrWSe��l���B��j;�ְ}M e[G9��Y��P���by�d�I�+����$/xjRk}np��ϐ��u�jJ�|��f7�\�Z7��}xdD]8���7�(9�� &����P3�������Gu����$��)��pG۽yb��
��ݗ����n-x�l��Gf�fW�z���l@���G��t�v�w�f�����D��0�>B¤`�v#���V��s���2Ou-W�n�����H͏�x�Y�IVs�-�5�w��j(7ܪ�<)���7������۽�A���i!�[ȇ��;m8�n��gP�:������  �Վ�ᵯ� ���?�C5,4�Gۓ� "�H���Y�ƫwu�g�,@�#�4r���^�����4Kě��ar�̻A���7{�1~	�b&��+D��ßZ�1%7�J�-�DH)�K�HVY��*�M�-���%$��/jS�k:�P�}"T�I�T������T�]��?����ښn �^�~M��*�=��y;1��?���X�	ɬ����lN���h�M��o펿�i�n�i��,�ݿ��~U�׿��(��`�X����'�0��?M�~�Y�&�O �t����E��1��^y_P�����*���,{��S����l�Վ�_"���\�ߗ��4�����Ӥ~A�o�����F<�}����2���������L����xt+v��U}���6k���f�����??M�����>�tM�I,�F�:v�n�a��`�i�����1谭Zo�[Y����f�d'�y)ү Ov^-R��.��4(��3��(�K�.wMeį���li�UM���V�=�v���;xp_廞dÆ0��3�ױ���l�t��2�6�����C�ƫB�^��ױP��v+e-�.i�b��N�.W3�Z�f5�ӱ����/�O�^�>X�0�ձ�+16B�UL����9x��L��ȣ����Y� �h@��u��)1GM���=F~�O\�h@�;F�:V_(�%�n�����Fh>�t��0
��B1֪�(�c�*F�Uw�w���%���=�]+P�k�N�#��V/v�Ϙ_uq#���nuN�V:T���A��e3�[�>����Z���$6/E�u��+:Mq"���3
�l�H��;�6qG�J���7����ے��o��#���<���*��		x�U���`@�K�՟���Vʙユ�*�Y9���xy��4��94]�[4�_���I��Xg�h�4�b��0-P![*�ZJk_x��S��&&�bȜ��^�[4�����.� L#-�/�A"�վRU�Zu1�ku�8r兏M�x���-V�^���F�KP�٩�B�j�cýV�А6/
\ǃ�Y��2�bA�"�������>�m��j�y���F�V��HuU"�ֈ��:�3���Xи(M�U�w�ގ��Z^:�5z�BJj�2*4p�1�Ʋ��@[�#أA���a��	����hgN�n�apX���ֆ���e-��ֺ�h��21q��e��ap���\je�B�w_<wG�pwF����;��B[5���҃^�m�E��_�
�2�V����qU!�51"~F�2#x����\�����J����e.�m��Z����*���Aw�e��i���Z���"���+��&>'��VÚ̵K�P��/��^�a�9��������m������̟.�Z�43�43b��������OU�ý��dq�u�-#Xè<wcO���s|�O��Z۩x��
��pKK��=�,�V�Rq$8p�����1��X�Hql�<���B����U[֑͌�����5G�4�DLp�<'��͑��v�FpG�p���F63&���݀)G5kݒy���l�w�v�d�3��h�ƋT��4\���Vz��厑�k���ϡ�:�jf�d�aU���0a��-�.2svWO� 4�wZxK�u,`T���B��@�������oՏ�\-һ���U��/��ŏ��Sz������/���?��{X-����ߕ��j�������PK   {c�X��_�  >  /   images/17d126d1-8a97-48c5-9cdb-beb53ba7b71c.png�XgPP���:�PZ�� �*"U@@z $*B���ބЃH/�� �{���ޔ�q3��~�����̾�y�;�����}1&F��@
<<<j]M�;�|�cd$w�Qs��!�ձB��qu������?��dCjY"�<G8������<N��.b>~�Y�J���!]Mu���=���v�/�����z[��l��։�Ll��BHJKu�9P��	�P~ۻw�����&2��D Xj���=í��¼�E��D���(���\��l�_4�(U�qOؿQ���;r�s������@u�$
��P��a׈~�KfJE��i���3���tL�OO~�����~��.L���(�,x�����Gy-�Ō�*��4�RϿ''�����42b�j�����-�<��v��ZJF��>4z��/��z�F�8\7d�&���>���ؼ�����		/���s���@<�fa#��	����09�z���ڵ�P��lI����a��>sO���72=1��SI�Y��'���哜i
~(�#Z�pG�<\���ssr��`�����B�)��(΅�����Hj��Rrޓx"S ��Y��]:��CΗE5�V���m-�"�ǵp���eD_Oh���\��V��B�����I"��u�X�i藻e#��D\�(�d�s�I1��]^Η�N��v�0�h8 )�37�+q�o�F�U��x��Z<��W0�\; d�ھ:�m�gN.�+��R=r�c����MZ �	��3Go1j�֩��}0Ä�"��h<\�IO�뱀�"[/��'G_�Oj�t��������u����J�s9�੣�2���]D{^������i|L�M��eW%��w�2�
���0O����߷�qZ[�B��,��@�Ǭ��ۺ�{mG�k,��0ZA����S~e���X��p��d��
]]y M��1^?Ν���e�e����:t�w��ۋ�5�ψJ7�N��՟юmB�A&%�$�4Z���Qe|$2 n���9�Wmw�����[��S���%�z~�9�T����#����W������ɽ{X3�p��1�j�I5}J�'�*���X�9��FFZ��ɓ��J�0ż|�̎��G� �^���j��O5^�z��iz^���Ky'k��bYJUю?�f9ϑu�����2$�busK��=(�|��n+��*�u�R���񎔀��w�_s�b��#d�?	\l.+��1IO5�ɶ�`OP�(��^��eM%,?�������=�i��b�(��P<kk����ż���`�	o/�Umqnŋ�_\�iq췪���b�yh���\���][;)�9S^T��k�J���$��jo�r#if�fNj��.��N*<� 7KK1�N��V�d���,�CZ�,�es�iDԷ���EV�~��C�s��3,�,x�Q4[a�mg�W���@IA
���Gޢ<��w����i'\}}�0_ϭ��?�p聈�R `�Ǐ���F�PPo~\�2�B����d�.�	�
|-���I�H˖C�)�wl�9��zwӼ��_Yy����c�ZsV�dn��530�dtv��8��"�:ZZ2�0��r34ig*p��&����e���3�Z�"0k5.�+���IР<-Н67]"��Ȗ����z�8m��eD���[� ZJ��F��y�>+=\3')�_�(�H�9:	�iɉ�18����"2����=
�t��G|�(lc�Ÿ���A�����s<��<����e��z��Ht>�MJ�!�-�CL$߱���G�;��vӰ}B�'���#�"jY_1��X$�ˈ��ω�U��Y֔�I#s�nAl�($J���ޣ��i!�#	Jm���h���j<�Kg�Tɮ^������������*0g�������'���_O��
�6�ҥ��i�>����5 �\վӏ��Kz��ZH4x�h~�s<!i�F$.��#w��;nO��h��4xG����^�o��a�����\�/��EDN�q����$��~QqE���4�&����⧳�RQ$�ҹ����\o�r)�P���4[.���HR���Ie�h�g����J����g1M�В�hK^Á�kG�7�����)s�������-=O�<Ɖ�^d\��.N���u�0�iݲ����`ε?�8��*1/�o�?A'�p��a���	�vV@���\}�$o��������K��\���B���`��ɐ2����ᗰ,�*�ow�u�uT�c�RA �M�e$�2yt�l4��Q�͏�~�>���R9���kU�^*��xλ(�;��z����vf)"㕫�g<�������ϟ������i�G��#�F.�%t;"����v��k5�EE$%$$�$�@��nS��f���e�M���ө�ѹ���gTvڒQ���=r�&Gt^�3��s(��ok��͆�R�Z��,�1���,���B�KYo����2����|L�l���U�[^��O^����
�����2`�Dy�0rQ*%��y�Fs�K�`v9��/��MLL����P��3������͛���)�v�P��)����>XCDȇ�P���i��'?:��z��Yu�����Vz;~\�D��1|��o�s�4�z����3'�D�Ga�/څ�g��~P)[v){��!ejjj_�GWf��ﲯsY���%�'��_hSnN��7�+���$�ak�
?����<l{#WG=<<b�Z���;�IgcY+�O�W������o|T������o\U�JG���pW�~{�Dbv-���F�	U-zf{�|a�/����+�3W�<Tm�p5Bm���-�[�F�Tra=8�/�%���}�nT��^4g�i�L�8���h7Br��)���B��ާ�ϷV�5 H�}��B���q�
���-Թhj��7Kv������
�S�^��	�!r�<Y�\ �֑ �\�x
++��Ly��ց:]-�8}��F�i�`Q�ilg��˲b�{k����>��C��>����%����2��k%�:�賋����V<mm��g�ƒ���J��h͒,��h��"4�� �P]�(������>�}�'>?���ٙ�J��	�o4˳���{�v� �rl8�A�$����-�,�]����(��T{�_�����NOK��ėj��p����3���]�d����fP'8���Mn����&��"#EoD`D��B�Q<"3���$[D��a��^�S��eïI�ES��y�����\x�Ѕ#����^�
���O�,Я��@&_ ���9z�G�-He��恔'���]Mm���JϪq��^�2�yJ8f��SI�+��XHN�PD�-=���o��v�"ڋL��I�A�c��JKu���0(~*��,[�G����
v�:�?�p*�T`��dwpz��o#���IM#D� �C��y��,G�A�b�QR��D�M�2��&J�����C�� �:�>jn����=T�DD���&kYiW��	d��AXe���k��`>o+ATO�_OTĳ�|�`��(�S�)6��$�1�T/aً�,��$��K�浨��X�e�L�j�é��x�[+���V�@��1���p=����&�S�B�z|�N��ږ�J�YL�?���J���!�A?)EV��+HLo\��'2�f]e�4(ZL�;��0�|�q$R0_���GN�9#Z���"?QGf�7ǉ�+�O�+D�o|�/Ҋ�W�N�p�2`�X��~ֹ�&�y3�U\��Ա+�w��D�6�-�!H���k�>��/��V���АK�۝-���j�J�>�Ւl����s��������ݷk}b�v]W<��}�يo�K��&�W֑�1 ��<����/��Q܆�=|�ID�a#<<��7ZL�1 üTFg�*��75�f��p7����5븥��a���˵����q�ڢkT�y�ۇ��M�-A�c���g�D1Ѥu?6=��ϱ���\��L<����ֲw��
,��l�G0�M�j��/��ޙO04��('}��F���h��j2�Fpǘ:X�L��'�]V��NN�%�&����	k0�&��u��}��wA�}��\{�����f�do�F��A�j�RbC�&5b3I���R	c���himݙ�hݩ/�A�,��S�X	F|`@��nH�3��_�L��2/۸��%����v[-�?�Zݟ�&zapj��$͘m�!{�M���l�������{�?�$;I�x�oh�.
u�7�!���Ѥ�b'|s�zg�-�e�H:`A�^����bk�u<�꟢1�,�볤�s�0�P���W����^��Pi91����_�g��m�X͎|8�}��L/x�(Ј�����A{w�~��5�N��Yv"w;���>e�(��Ũ|6�h��(`	��W��s��|z"Q&$��|I�CqR#���W��C�cYcھpw־�ϛ����O&o�٫���k�k����7ׂ�c������F�}_�<J|6n�ls�C|�hW���e�]�	TT���$-�!�3+�r�ez�8��8�3��ۙ����7��c����'�ܞ��� BP��;2d`�	����<�Y��8U��vt�n!���#I.���I�u��H(ueY{��k#�X��|�5�9|��y����P��>
G�U1"�E6��Y7�~�IP�� lBy6'�T�m��Ҹ�}&^�BD
��#�d�_p4	��{��� �>۔�o��렡��������+C7��س�?�q�/�O<K&ʷ�	�)����*;�.�q�aD�ב���~�K����q�o�rF�Nܣ�Vsx��XH��������?�����`�s��%]�~t�U�y#�磪Q�Fn��!A����!�x��=�)ɛ��dee���2�9�+ �����W��'�fzqV�.��j_:�6�Cɜ�&�[n3ע<�S�P��d;�0+v�M֥��9��>?�8Ra�TЎc\�����M�3��vH(	�������dy�>��R�u#��&Ʊ���F�8���%�t����l�^6;�4C�@�-�^A�4�����?`0�XY��ʡ~����@~Cߔ7[b:��գϻY4�{����+��{w�Xgz��D� �x��K��������^��h\�[QCC�a����0���sħ,ߌ:��h!>�^��:6��"��*�,1�<��P9�.951Q�iiiѥ��i�X�ǙW�y�I��>-��g��nJ=��Z�����t����AX��W<�kA��*����l=���� �	4�ި!�$^�3'E>zN���MP{Eu{&�����ґ�_l�ߓ�����,���b���E��|����$i? qU��H�[�#��z���'�'��U� ��n�T��rx��l�O2EmV�SQk�$)�����A�~7����Q[i{�U�0��&��5ʖ+`�S�遇���ۨ�6��ɎZ����Uq�
W۪��N�PN3��'�8��I��������)�>[�x��*ب��i�}�V�vK�5�qM��{cr��Ud ��)�^끕^�'��i'b�ӥ�� ]J�F$�tn���o�t���b'�.��Ï��%1���c"�O�K:�J�/�<��o �� ��\-^2�7��)���%�Ա.K��ՓW������*j;����m=�N�jGI$ɇ�tY��uf�J:�(V���*��'�b&�̈́�s�NN$e��9[e��J��R,=2e7��lË�T��T}��N��U��>i5�1+��W�X��Zu˿�\���ն��"�c?
Oq���^�|n�~qz�؁�ӛUUu�0/�Ԭ�``=G�#_u��E�֝AZk���8�&�O�6L�a5��'��%R#����s�;�8Vx�-�%��V�J������V8��i'���ȹ!�*S}�`�1�WM<|r�9~����rTYq��A�,q8��j1�G@p���W�;��o /�4C^�����8;p�!���W���C�Oo�REӵ�}ձx[�o�LI��;U��ə7ޜ�.�f?�C����Ozi4>����>�.�XhL��|���V�n�nWf�l6���Ǐ��ӈ�#���z(�ǚtݝ��E�E
IYeq.DYC*��F50婻b:22t��ITi[K�t�ƹ�}�tFdYt��j�"<j�g��#���5U��}6����ӂGR��τ�����ʭNx'�,��.���$F�tV4���Ә2h17�D�Q��ΑY������t~���������-�A�{�x���u���T��q7��S��ˢ���t�����W
0Ƃlf�G:���/Z*x�:�!��_^��\�u�I�)��{���� <�;�"�lɺd3��$�"��>zf0<:�+�]���<ARwPDR��&�$�l�����OHiD�o<���xw��e���8��PK   )_�X�C��z �� /   images/182aae98-c01f-41d5-bd55-0eb3a1cf7144.png|�eXU]��(��.�N�A@6�JH7�H�t�:)���n��ݍ�t7�������9׹���{�k�1�q�s-B^�(����@��T�Ah�ʆu\��q ���\ ��<����=�H�*���h��a������v�u13u2�u|c��+IAL�S���g�v��/y��_��y����PQ>~�'U�]zu��i���;�#ߐ�ʂ��!�Y�Os%�l|���1�Џ�(��7���>�So.S\N۽����o�KJ����?�H1���-9����OJ��v��^JR�e3��P��P[$�d��Պ5�F*�� <"@U��H}��:�d��E��XPF���?aF#���^6��1T�b�Z�����y���!3w��+��B|������-�S���E'$�p�մ��չ32JKO������ק���Ӭ���
���g��4t�Ɋ��c���ț���		Q�����)faem�WE��
n��������a���w�*�Ǐ�?�W��:��,/���Ζ��uH��&/��`Н�<�igZ(~�a���������ז�+��N�3w��񰱱�������������T���E}��s��s�!k4��Kɻ��<��-�0K����[j�}�5�|�,?Y��M���BLE�Ar�zqq��G^>�O���r��`�1�Du=���c��kku�Fs�������-�'~x��:��7��nnn�Z���A����!%6�	IW\O���]�}^�����Y�ҤrO15uHI	�B~F���<L_�[���xa�J��l�D}Û�����|�tbﻻ��m�AGg��������Ȏ�q�e�������޿G�DV�|�k�F��{z����=��͵�����Zh��r���Ar�ěN�]I+����}{;LSS��Z������������W����^�U��K&�	����<kk��^�1��@|&��pHk�3���O��o�$�����wc����-��Lw���+*4�ꛚ�6FsI��x)5��2����y�����DddyF�ppq�45?>����O�3���?Y"=/�{����Gܳ���c�oF���w��O���^]�mh�����>���"�̌r�g��9��f66����:cE�w
������2k��u?�
4��H��#Tpk��EͶ����V~�y�$��8�ٚR���
k��w��X��|��=
J���Bwf����2�?:���5�$}�^ԣS	OĘ�G��@�̎ w����ETT��_��質��M���T?I�Y>Ub*Wa=�(\}�� _el����$�?|�*e>��R�ڞB5�ۙ��p��^P5���_�P��E�^�/1����/��U�M�	0FA������n�����SO/�Ʒ���Ab�X߯@�=1�wJ'CLJ"��Xz�>�Gx ܡI�ſ�T��EC��k��x����6Z�)D�6!��!.(����̧H���D�b;;������mc;��)�}�|����8	7�ްs?�(��?����#'�V�B���g�8c���͚��j-x(:�fP�Ү�^:�"�D�:j����ڽ��ڃ)d��`�0K���̧��[��v��y�2D)���|ԓpE���8��D��;,���Ѱ��g�1�4���'J�1br"\`�^��@�qMe���%2�g�=������QpZ�(pY��P����Hg1�������xvp0<ङa+�Я�d�Ǡ#���v����IU������2A��t'�_���{�QZL!3���/G�
���yDP0����G�nL��b�O�`�=gޗ�H3d�Nw�X�1���$먧q ���$�NrW�F��z�+rٌ�?5j�9���g�A�X�P!�k^h�[��'��)#D��z'5y:|��J-	����h�~y9����x���(L�U$���#�ƖUW�����m*�ʧ !%���ʰ�M�W��c�������C�ٳ2�������n�T�&�R�heL|f��D��n�<�I���6Dh�����y_��Y$���V
��� ĵ0�����gX1�%[sc���y�Ijd���H�PT�9����V�&�ԧXG�{���b����8Q,��=N�Yd1"�G��EE�N��۬�n]��0���F���b����S�3M\ ��&�u}��b��ID�2�����%�}%ݜa���OX��l����QJ~��F[�Ӊ;�o��+�aF�c9�QA!����P�'C�j@�h5��S�0���D3�;��������y��7���cd��%�������p�q��׷��1,�2Oy檅��������ҧ2KF���I-AI2�+��E^!�xiiic��\M�+Z���,�� ��e�D�>/�|e�S�w)I�Y.p�i����cOϚ��4( �+8�"=���x�����eG�Y,��(R���y���EP����w��D�NBL��ht�ۅ_�����'�={FDB��œ�칒��Vm����� �۶N�������YY�Yw)�h]�����C��J�ݖ��_���>�Wt888���y��K[[��>G/��6��5�5^8uV��KN^�L^���o�.�/+��8��Y��
j�I�n!��\��\?O�/���3^~�hp :�7��>^�����s�T	�+A�4]l�~1�4Ӷ����V�Jb�EN���b��P_,�>��(		�2
-%�p�~�4�$:�)��x���#������B��-��pc��,��	2�**Ex��p߲�B�x/C
�ٯE�՝@�S�y�́o��Q6z����|EY4��A�uC1h�m�B�����������p�A�(���w
�SO��J)c�߅��*:�1�Ͷ�f;0uq�I:�2�5T���'�� (+�t�ĉ���� ��`��[���2yF�(���Ѐ�(K�E
�N�$�������DǋJq�&B[�A�z�tk༌�������`�S�s��m��%��ĸK��ъ��5�[�����;����1?��P~hs�y�I7�xQ'�%�Cݿ��*>�:M$�裝c��?��������ϡ���BM%��_��m�>X�� 
/�D�����%�Ei�=|�x ���1Q�9!#-u]p|�Ϳ�>E����f.�B-s�R��A>Ә0F�F�P�s3C��]�%�F�z�:��&���Wѵ�hjZ�%��8�W=Zi�5���Az���99y�T/��+�c�Լ���ׯ����w0Hˣa�p�����aڇ]5ޣ���s`�j�I
��m�ыLK��Q8��c��]
}G4�Z�J�*,���5������4\�B[�
��N���ڂ����k�����`��c�.�/ɐ8����E������3�F[w|O�x�`-�B�4o����&�S�w�u#N��v&l��ޣV�][��g���~�JW*��"�c>˔駄�����?�<�J
��������@fe:'�L���8��?�7pI�n��-&�3gøT端���זR"�]��}�f���X�!h�q@�1�Uv�h�~d��Pl�1���>���ī��P�b��F(��̙V��CD��Nh�q!ΐx�諯}l[��n{�{�c\
*m昦m�;E���(�'-w���$�����"N��F�$��	������\g�Ej�]�!&ѡS��Q�/D����2	�;O��m��BPM� ��/*"[�"2��^R)��tJ��7���C��A�wj�%%>�e��	|���_`�!T]?Ψt�T�*4Ę��h�:C6XY�ԧ�Vi�b�����ɠ!�g�d�V�=8��j�|	}��F�uZ�c��J)km��C�Wկ�ape��t�)��4>��>!��8��K뼡n!b�$$�s�[|lu����� �HD���F.g����R%Q	u�����'@�����1y!ϟFϿۿV�<����R"t���A\��M�yh͡8"���g��0RH��o������zdzqd���!6� ���d��-U�+�c[��~�:��=�w�MM%j_�f�H��~��g^cJ�>������Q��}���i�\�3V�9񉆬�N���:~C��a����|>�:D��~2����P���JS��ڪ;*��p���n��<������B�!k*���*YF��v�}b�=�Dj��	�#W��"`��7�-X�l���>P���&1�.p�T���AV�y��a�?Ň�gv��}�mu��/�ܾ��L�2Ě��+�b��� ��d��-U.�����ՂX�,�h��4����,PCo��m�S���mW~�%7γ���gB�Zޕ�?��1yG��zc���5*��O�w��m����\M';�Y�~
g^����	��|Nf�㙽�M[ٚ���Z=�E�H���CM�ܛÊM�s����c4Ŗ��?..����z���ʦ@���P�=�� ��	NG��,��a��_�a��٤K�0�h�*�Ϝ�j�Ԉ���U���S�a%|��H��NO�����'BY/� �����{Ľm�癟ڋ?si�60�:��~�Z�b����j���#� !��<�,d�ǽo�=~�q�eμ�?˾߉��dK����M3r�����^jX߄�hBhV�es�����l!D�K\_�r޿�E��0QL/E�c9��=89�h�F�b:���V�H�y�:u��2�f�o�7$B�=ŉ9��{lh��e��RD�v����%����/�}BC��-Nl#�,G�l9�Q�܆��!ۤ����2߲G~�7��{	T�Z0z��ʒ�x���1�x�w�D(+�_�eV� �ǝ$`�P���*����U�C>�����V����S;I�Ho~A���h�i�"V{�TA���GM;kzq_�E�8N�PF��C��6�Rez���G�C'�W[[���1��#%�GMMM&!!r-�y)���#vn�cW�$		�x>�S�1�� /[%����W��L���xrv�2���^��M]v�YGG��۟�/��$Iz�dff���j־�q�GΙ��
��'�9���
Kkz�s�8/�b�������>���տ�`T0CVsǓNr|�f���i8�>sB�n��ҳ �A���_g��)쮟�̈�oS{Kcacc��|�Cޞ��x2�gc8�����y�e?Ӄ�EFr�^���%��UuwVI��������/����"�|}3$�lhYZCHٜ�֔���<6����YxC��8LDK��D6���,�%:ZMO/[��.�����q�������(*&���˽����������s,�ZAC*8�\Vy���ǩ����5n����������DjN�ӧO������G���.��//�S1���=�p�TAU��s���X�h��Q_�@4�1�@�k��I::Uq��CD��,Ы�V�V����;�������+��{/X�%g?J���a$SH�(��t�m�J���P��HO���c�
�f�a�v���JĎ?5���*�roޔMDd$�/x����_����a���h�Ap
�e�����Q����bfO{OO��W���T<i�;�������(�&��#��fR�����Ғ=�g?F�ӌī"�DE�K�o�3�#0`�~4o�#fໝ�$B3��Z9<�(��=��Ys�dd�G���)sS�	sR�z癆���7�уD�]m߷���~2��)V�m��H$]GEv� _.S���O���D9�������W���YƢ��	0�x�'S�(ez���j��ב+�m�U��*-+���U������g��·����4��ލ���p�r���l�������Hd�G9ly(m����Q9��1�p���e���sh8mLeS���Y|*��
�Oq�x�߷��E��u^Zie�p�W��S铁E�TS*�����_�	�YG�����΅�5h���'�C�������;�%Sv�Ј�̳z6z��*:��JON�������R��vh��F������k�ږe���P�C�(��E���L���.��a����M��w��ձ.����d���h�p��(���N_D���*!!o��0�&DV�9؏�Ã�������t�9=��Q�� ��2��k����r�W0�#o�x�g� +%-'��ٙ7#jw���\�^�6��߿I�A�z�r	�z�x�|a��M�l]l�a��9��f�zk��eU��}�'����+Vݜ�[5Ե�ɕ$��		�e�M VyX����l�:��˽	@���|^��A��ΖĪuTQ���
Ł��Ρt�d�է�nD)�53���������/�B;�n�8�er8Y�̄�Ȥ�G��41
��5oVCg��Q[IY�vrkRH6mp�T�������g�d�wò������Z8�nz�M5�U�c6�Nٰ��q�]�*Z{S�H�v���Z�/��O�d:~ja���8�G�<�jd&�ci�NI��h�B7�1���>�G�򪭆���W��P�bc���3���J4�����D�
�5+���Rk�|[��KL`ٟ��dkB��:���M�y�N��%S6�>�u�<ݧ�����A> �Q�r�e
>H���7�N�n��������-�A4��Yˏ�"XP͸Zd!��3fb���u1�
0�}�c�d�H�p��u׏���xo��./��	^�M3cY�;;1=*�#{l8�������WZz,N.�cl�O���'�͓�V��[�:�^B��X�x\<[��{i�)u�\��;��y|l���a�XA�Ƿt�f1�(�_������~���Z�GVL��π-T�)w��U�*{�yz�i���//Eg���}�k�dMY�Q���*��7I���$)�X��:�"h�����2�o�n3�"�ޜz�>k�{,}Ьڴ~����	��B��n���$Ì�Jƶr������5��t�/��Ma�/�rfsC�]��ة,>�r�{s�_N�����,���I4-R᥺����ڵ2=VM�4ք#�W0w������{>�_���
�x�O#åC��y"
��;G�y����j�8�c-PTga��������/(���~_%)�j�~���d¤��vbT�������EF0yyfnn<�u]�ݏ��i899�V>�01���3KK�P�Vڌ	����$�X^K01A?~�H���U�E��ԄEHH���ǧ��i��{L�Q}��������?��4�D�A5����3�%��͙<Y��\ZZ*��<:<L����/�10��V����ҽ23#&'�`y��M�OHw�����[,\\�d��^��~�7F�~��O�ӎ��8����ۙ��)�i���@e��·�����sƏ���s˔���Imh�-�ky�eff����w~u�
H%�JQ����ٙB��)���l�. �P�4��*���@|Z��ŭ�0Z���Rv!Z����&5N�����O�����O���C$��q���[�|A>�Z^YA.{�$--0�6�;N[�<�1�/�J��xA�_eg�+��B�0߀|P=����>�*��"*JU�0��{/^�x)Yq�OKc	�n�! x�?[�ܶ������k�c{���h���� "��� lȒ���J`VV�$$$/���Fs5:�����M��i�����E� �WR2����u�Ǭ�7� �#�#�F��$�f��*�/d`�vB��X�7mC���H�-8�(~/��44R�V�z�eSᒴ(�<U����1�&i��[����'��p:(c9
sQ��}5=4�ڥyq��L������<i�S;���I�  W��D�ݸc�ˍ�
�
N..�{Ϟ?�����쌲èɷ��x�����OLyS
>c��Y����`v>�O��52�:�Y��ן_�zջ����b�CFA1<��c=��|���]�׷�c!S.�����~���\���E��ͥ�
 �_{��=x��|���D+���[W�A�����ֻ�����?}�4�
Ro�������w!�X@�a��Hz[a���F�PrWd|�OWX�����f�F}���k���P��J�Z���mRg�r��/9���x�2'�v8�PPP\�ϝ����27��F�U㴄Z�W�����3 ��`����rGXhPo��&�?�=�MG�#���S��&oo��MA�KI%k>MW����aU�1Y���]�{�am�U~EE��Ձ$�OsY{!+�����<��B����V���r�WW__��z��c��V����=@fX���$$�Z�gd|��>P(on�,.:�� �0w^�ٓ�(�nLy��	���x�}�S�$��9�<&!�Cm�ap'�~W���m�...,FR�|y���"����J�Ao[�F�بL���ֶ��5f^�H�GJ@ ���X�}���қ�߭�HQ��A�_����_n��{���	jkLb�s@Q�Oчș���C�WP�Y�������V�v���Ҩ�+���\0�(���B��Ę�F9������v;�
 �$}�B�_���1�H7cm޿�[|�,GV*'�I���=�;�� �+�+��������h�sʄ�&���־d���c�Է�X|��J�nw��(��W� �CӍ>��.$켼Yҷ�潷xp��\9砍��Oi�Hz�����)�f��~J3����*�+D��0���*��lƯUI%���r�Pq�I��C�c��$f}̙�����HFLL,m��Y���Ç1q�z�O�nt�����=zvW�e�Ս�U@x��T���s�k��^�5tn�c�����@\
vDu%���t[��lmyZ2��n�����_z��eu"��gǛ#��ҭ�/��;�oD�WV�0+˩��"�pG���8&�M�6�83cbc�&K��%|	�# d|�q�+�R����RT�|�j��ښ��lާ�*z���G%���d�u\�u$�ɑHv,�<��/<��ə�3�k٤����a��jq�mw��;��[�@<�^��*{�2��|[�J���WWՂ跋F2�/�����O�^/4 ��\w�q�$�������CR���Z��ηGz`!2�-ѽ�SP��o�x��3@V����$���S�UX��O����~�:#g$-/�{j��S�x,b� �UC%I��$AOb�bcuu�u����n��;c�E�a�m�:ď��*�F�H�� ^� �H�J
ajz6�O��2�������?�~ۥ�/��V888D��B��{Mm������"�������|��e������?�si���<�3�4ֽO�C�V���
"��;����}+FFF<��X>�ۥ�[ �ܕ�0�F��}�+�0]n9?�d4�k�#Ta�����c���s�GPAW�Õ���d�5飫��_�(��Ɍ��S|����uZ i�k�������˥C�B����yˏ$���Sj3�Yn�%�i�E��#z�,�����r�1 �no8�հ�{l��ݻw_Z��d`���*Ը�s���`5��՟����f����2���k���v��
쓭��A�7Wgf`7���f�$�ջ�	��HMe�X�G�j_`nQ����C�Da|�.�F��ԏ.�]��?��Yx9^�gі�ȏ&������h�}{�/%���"P���h��gY�t�Cʦ��M���Jm,�2%�����|)�qT�D|��vln�"�X��&��ڂÊ �ӂ2"L+-&F������_ �9�h,Ws��(�m�Ҏ۸����u��B$��������<�}�;xû��d�_bO4���9�t߁�S='^��z}q$���6�@l5����ރGf�pY�K�E^ꢖ��YY���8��kb�vZzv��Q�F�zu^a�ɗ�3:q*( $�[q�\�SG6?��g�j5�2�}�瀊���������<�������B����VD/K����"9�b*���.�{I�c����F�q)ѱ)�JE���v��ʒ���`~�,V=���l�FB%<v�T�NȤ�?��D�F
#F�qZ�eg$�pD*)1��X��� ��:;�{�Fv�+�M��6G��Ϩ���"]ѥ baaa���SE��g�؋�=�F�!��6�%�(�#�t��pɊX���(��F����G9���i�b5]�f4d�|�E�e⾾�ؓ��|�O�xԏ�%���MYed'<�FB�N�L��mEKeE���d	bbbM�
6#Y��H#�����A 7�'�[Q����Z_A����� �B��d	���J{�*U�����$[%��� [�]���M���������M�����R�����'��t��X�j�TM�� i��{���8|q�n�E%d���|{�<F]i?���ֺ�/���[����
�FЊd��А�u�\�9�<��������y�+��U���g�������81WZ=v���T��|�Z���-`@�)Q���z�����niQ�
���T�/�]*��X��#O�Β�w�17E��&*�@i�yN���1���M��� �R/O�4 �ټ9[�oԁ��Β�T<=k����\�zoo��'�{.cO7x=���k,��M�1�u�Y�n��W U�DFJ*���Ӈ�T���qS^ �a�,���
.�f�:pԮ%�nM�C����S}��$�hl9��V��Ѐ��3vs:ٞ�x�����5K��ʊ\��=I�I�M�Ա��d�b!���B�n��n��:������?Nڗ�F#��"��=i�u�ptt4y�����8'��ۓ1�U��ocVf},z��eU���+e�	7�P�<`���{}Ga0`E^�Mp�	�����o�w*�3���cB�UF�Ÿ;8�v���ly����9�@r��Q
��(;�M��oLb�x�`Ttb"�-�S䫤Suˀ#���!�,���t�k:OHjD�9\v���1ȫ�Rhh(lK%��)���yM9 ��8AR�s��~�;�_�f��v����C�k��x�I�Al��}	P"7�4S�?�ӷh[X0�����.(z�KUM젲l&v=�7�'�x��P7���Υ�U�����L�|�x����?.���s+�Ȼ���Ks���Ms��a%�|����`&7#�����`%TcО�|k�8> W+?�`e�B(g�����Y�r\LLWk��۫���n������j��cS*k��� �QVg�9����2!ȅa��aK���ܗ���2�"3��������Tw
Y�v{{{��,uˠ�U�͙�,���ny�J��t@��Z/�`v�1�V��]��,M/����Tl�;H"� ua�@]��l����V� �-����U?9�����H���^`�a���"�$�~�����U��r��;^��<z��o2�1��p׉Yːr�C6(�=F�A��5��(TW!b>���#A�Ъ�0]_)`e�����x�k.j_A���-�~�֗&z�<�ٞo���#��^,wX���,�R������~a�F���{�ۖ��_6�$+��2)@lMSeY�r@��)�]�>�u �*+k�gg'����k�N�l���VS�YX�<����F�3d1Ns��ACCC���BV���}����D���1*���h�i�P�;�r��z������o;ee�x���7E>�Լ�sA���b载���M���(���]�W ���e*\�XXP?Iw5�exuuu �\�uu���j@�����4Y̌7.�1h�IKcA���Ix��O}���BZ$���5������OҼӫ?����e~,a@V�9QV��.�WW�o�ަ�pi�\̣a��4���I&.4����'�}�� 2�����l��3Œ�3�:yvd��2~��x;�P2::��ֆ7��S|���T����k�օ����V���#ȃ��ә4��9����>.n�ˀ��e7(-����d�R��g>�_�X�Dx@�(���˽���B��J)�S�g�4@�i�Є��܊����=�茻R�_z�x�j?SE����:K\��!ZI�@��%>��py�I�_Fg��2�p~�M��
��b���KeV���X���t���i?�-Wa��n\
n�sP�a��T�B��P몪�\��E(+)����Ңc�⫠˚�kKK4�����j�Ik|5H��u�4����Yb�G3T��Dn���рY��n�+�d0�-��6u��$`�-�fȟs�4{��q�����V����gۢoK����
}����7Vvv���������{�̞{^�ut�}o�G�Җ�I8�����A�z���o@�P��p�PSS�z�n$�{}��LdA�ƆӢ���yo��'ȭA>[���o#Ș����f'U��"�5^8��ʈ|�%�3%�mw��*T���kh8��R�eJ~���%�ׯ"���&�z{�$OF5 <��ބ�R>USW��.k�?�s~�����t��O����\��&��C"b�wb.k�`�[?����G��SJ'���I]��K���s+$�/����d}`I� �n��XOO�s�&D�$@z_��s0�˗�.�OLĀ���86GH���<�3VV��m
�";//E2b�܆�����t�ߥE�hkS�6]9@�]C�
f=q<e�Fu��b�Վ��I�N�<H���=����=�J9���T���Q�롵��o#gg���.�3c����y�s�r�]�����/6br�{�;%A�!���� �TGH[қ;H��c�*'/�2+�'C���Sp	qՓ�����YA��*����%T)�@i�ȵ�c��q��I�ˁD��BSHTq�f�yO4p4�*���"�$�X�~�o�+�kpW�J�*٤ZM+���w���ՙYn�kg"����=£��k<&٭]g0S�Y�p�x���!jn���p�����t�q��@d���vb�k�ɬc���[P,i,������qD�Fb����[�k	))z�b���z�j�x<�#��w??`��}���)|վvu)-�W�ӕ����	��Fx��YY��S�z/K�zj��\��JD�ԗ�����ි�J2�0\XQ�����.x5Yb�1Q���'С@�ִ=���%��e�;4�P��쭣���J�E|�*]8ٚ�R���e���W�F6�;
ڝ��N����[��d@������a���U�m��3J{��LQLP�H��B�>ۍ��w2�V}t����o#�����q �r�#��-��<|q223C�	����齆�$�����g>�9ֈ�f�����[l=��*с��U_�$�(2_�DfBږN����{
	�t���/$�.v����9�~P� ��z-Õ-�k�C_�㣕��Tυ�	�C�%	�?I���m�}~��=1c�7oU�?���R��o�7j��_�<�w	���`��E���ϣ�c�`A����h-�؄�WLN�NmĔ=MAs��%T��4�Iȁ�-5�$ʾ�����H���Cd� ��*'�]j�qr�$3g,{�R�5���X�O�5����|����|	se��!l��oc���򗧻s��䔾a���~zt�e����`�'�/dN���)"�����뛈c�Ǐ�F�㞏������LYg���.hz0[벾����ܼl?!!᫘�}�s���fQQ*@H��>��cU��u��.�����3R�p�ud�?�I�2�;�O��p_`��_߆�}d���8\7!���� �v�W�[.��|�&����Ԇ����K��_K&!��ďD5���G[�A��"O~��"&%e����t�D����%%5��p��0�C�cPPX馫x�
t$xma����)�:M�&6j��={�IsSN3!ȋj�bY��R��>��[q�� ���r�Wqy���qV�1������y�0z<)��1+xdf���Wj��H�N����x)^�0�,��U@L2@ ��	үW�E��lB4�UBh�l_��/�g��H�����C6��� ���,�����9F�J�{�Wk}�SF�-��U�o~+�#���C �|9]a��..���rl:���g\ZZ��qf5�;�Z�ݙ�N�؛.L�����&�o�cӻ�b>�׶>cO��fk~P!٪��	9(��v/@�
��]]|I��b_�S��>�?6����=��D�G�O!{���h��ځH���3�y{��s�>:OM˩ư���|��-�p� J�p^F�>ݶv�j���ﮨs���B �Mw�,��tgF����߫��㒿WW�	tṔ`�"kc�w�mh��Q�$,dbb��jB�[��@�]��ZT�T�1S�üW����B>���4��=&x�8o�|<㼂�Vx���x���u�f�SEEŒoA,�����/:�R7�n�[����>Oe�J")�� �P���l��k��9H �Da�d��!��~��?�NK	��"�ľs}w��Gޟ�6:P�Iy0|��f�ۮ*[n���#///<���E�v'�Qz>KA��u�"�4`vXXX-�s�?���X���o�����<��h-4h�P�9��N+*)�ֱ��C/%��x�zW˓��ޅ��BtpSD���n�OC��
�>�H�9�u�%.����U�����缼�pc���rs��XI}�S�xDqQ�������s�av�'��_�%~�ʎS�ِ[.�.&�'������hv���r=��٩an^n��ACZ`���P8��r�VO����[�����|�p_�L\J^݆j)�Y垊ѣk��������Xܪ̔L|��RU��̀�kij�pp(�����ڷ��/���?K���Z�;��å$#��c����<d�Ovߙ�2.AH����NUy:Sng��>I��pZY�T��#��v�>�Q!�\��1		8f�����v�c3��H�o@.�����F��]���.4�vHި�1�E�pW���l]�  y,������I&����&�)?� S���Wn�ᝋ^������g�4�C ���S����y���	�}~hOQ���������������B���{�6m럹@0�l�����k�d�ӐQR�zo��p� (�X���E�����6**���B>�#��_�ձ�/���W���g�L���u�Sj2���V��<�8D�<��uԨ��J����
�#OA.�l�t9�T�)��f�{�~�F�GnO�'˷;�Q�3OxZ�Eoq��h��g@p�S���Eu
8}`�=�P�^����C�
�# t������Hz��


aYe���R?��1K�n|��	�k�V�|��h�P<3�
pn�*�љ����	33�n�U���;����}�w�[��"Z���wr����	Z:�(%�x�MWه�
��S� �m_�YXX�Mvf��l�s�J*��XX0�Ҕ/la&\��@�=:��|���@�>+K�ۖv���D�t�w����3��:��j*U�ۨN��! �@�f���>tߝi�@B������ BF��ˆ�~�(��9ggg��W�F��'��_��!����bx���}ΪjZ��hi�.��(v�x������3��Me�OMM�%h�&���鯱���dUX=�����L�����שee�*�ҁ�����	�e
j���	�w����t`j[Q��ii�(iL����v��a.Pҿ��.#p���w����L��ȉoV�05uP1w�)����?ܶ��^�״�pK�ӊ�����s�����/\��7Y�߱�V�ud��V�as$���W����F���!h��2�fvlfv�f�Kx��Tf�aT�;/���lӱ>�����3~���4O
3n�/(��9J9
��7�gB[��
%��Q�q���P�;��x�Ļ���x,-/h%eF_��J߬>k8��I���?)P���ЩgVV9a!!�g�s���V�ޓ�׶�l+H(2�����,�m�Eߛn�*����0Y��:��!Ec�&&kS��".m��@3��'`����������.'o�zd������!�չ�h���]i-�88���66�f=���]s��W2�F'��X��
�H��q�F@�q�[���W���%D?�..�D(�m�_�qn�%H ������6�&a����VϬ���JA��Gto��k
�;aC�O�Ɔ�Z��h��]0�4�<�'�F�ܯϝf����l EJ�j�)A��*�WŠO6x�[)�¾?������@}jj������'3 x�=|�{�j5w��_�`s��m3���� ���y̨XZs��a�K��t�d{MO�i�ݚ!X��Ef��c//1a�I���Í>S�����su�HHI� ��<��9����)*B���O�d�;&vߞd���2C>&�)���{vW<-=��y�I�(�64�%���˯EӀ5B�А���X���O~ڡ��^��&d� Nu��#�8��VV̒ny^hk�'A86�0�`��`%�YT��ښsܿ9�ё�
"y�r��`R��QP�T���?H��k���鏹d�r�m�`{��>;�U[��s��9��y:���}G���:m��az7C!��;?�,;��f{R ї�3P�
�~�u��N
ŷ���	#phO�tR�K�1�Y�D��#����tN�����+!f{%��.L'�@k����Lz�ڠ-���~1���=$��$%/;�W��y@�T���B��>g�o~c���M�w��d�qf�X?�!�,�=��?x�&K�]�ܘW!��:�Y��x;����b����Xv�%mxX]�s��Ǡ*|�7A�V�������(235f���� ׋����%]��	Y�ga��.*��4y�����&���n��w�4�����j4����~ ��Ӈ�JKK���9v���<8�X}^xGBV��iNUܪ�U�����������}�j(-��6Z�G��R+�%�{r��F��Z�;c:&n�XY.�����ic���*D��������VV�Ib~W�z^��~E)�ǂ��������4M�[퉷����Pz0M>l�(AZ�*;�d��~�{Y���&�_n�!_����e���[��D�c�fll��v,=��d	X�`����o�<���t[*�1d���Y{��R� }���%�ďUY]�踸'��ȷ��o�AZ\
n������� �ji�=RR������n�.�C�S@D��DD��Ni��.�����~���Aϳq��̼��ϼ3{�6����J��E��m�,Q�绯fN=@G�hjj�(�����p�'-1nɀ����f������(~B̍��U��;�Z\�̙:�]��mi��,;Z�Gc�Q�7(�g^Q
�ys�gy�]#ystSV0���7�C�9I�����·*�%slv*��g>��Dت������6�!�;NUO/2�E�y�яru�vp��T>3\sl�����4��r�a4+�LQ�B-yeeL��CɁT�a&����$^;bh.�+��Ԩ�RE���i��HH���/	�p�Wcĺ���=L�ؑ -�Ï;LT��O\<��E~y##��
�TmflRR�XS0LS%���ښ�@�2I�R��\ӵ�JO�V˕)jV���,��gX͍�7I�ɩr8if�ύ�/���gfw�fppqq-0;###���.t����?��'H����/��#Y�Qb?߰9SYh�U�Z걕�H����qk��v�����nv �z��������4*�^*(t�dK�[�W����>�Js^{�Ā���E����ԯh�C ��g�A�|�qh2��Z]��*��^����L�E}��q1S ^+N hu�TZ��4���S���3�'/�<����C�YdM�ڠ���a��ݭ�:���GMJY.���6V9��i��e�m��FdT��F�����w՛)ʅ�]���\^�]�n �@UQ����R�	`�W��ݑ ����cbD��jjR�##�f\�����TU���v�A����RΜ������U��>����\����t	��s�Y���k�s 4t+,P�N7A&{5��Cm;���n����H���-ׯ_���۳M�����W���i�l�Xu/3K��s%�NA+
�_���<�W����Z�]���ϯ�����U��<��Bk;�\��a�	�EY��[n:�����~�K5��rL�="c����7P��Ƿo055yy�X`��G@�wnO^?-�0�H/7�C��B��6m��J'���Նn�k���Ȗk��P7�W���G�����7�'&z���ǡ��rXl�,o@G��O��yO��CK����k:0p��[�w���

��}u[�~����} �����oL\JNI���u?T9ԋx�Jlll��A������6�v�Q4�R^`��JK#�
���:����;�{_�w(�(�����^��Epuu��ꉡ�q�}���c�c&LX���P	;�)@K� ���9���,l��Gd��B[P��a��u�ٿ��JHH@S�#%�|3Y��@�_���S7W�՗��cg�R��;99j�A���E����)�V��)�J�Zs��/۠�"��T!�S���v5^��	�Dv[�kB�����g����I!��ܹ�$�$� T�'8�X;��t�|���s����c�]�?�����s�8Z����'��=ʇr���'<��S�'qe��ۆ��^��0�����L���rb!�F?�Ǟ��h��A�=R!���6������?~�QTĀG@ i<8����,���&~NN6>>b�r8�����y-F?�P��d_�z]�����=`h)Yَ�E
�tLB6�F秠w�GF��ϖ76���9J��2B���m��$���oJy5AoAd���&���ЏD�q�V'��?�G�"X�N���Ԙt��}������g�:�V$��=��8 ��/��|��?���'K���}��}�+`� �].yl&�8x����#dM�M�Ͻ��eL�>>�^�%�v<� Ԕ��򦶇�������5+99����^��v����%E�֣�o:�"�:u42pҽ=��K+<2	�F����&wP�1����N�?G���o�����o:�`Np� �����C�����щ/���c/��'+���~��ĩ�R�al���U�r��=����~���'\�ǡ�Y���/q��v;?�y��Ӿ�o;>��g1��[(%,%���N���٩�H������|���N!zuۙ4��DI���~>=b�3e�Q��Z����'ay����V�E���N�܇$+:�[�R���;K������P��ow����f������E����Oel�Ҩ�q���x�=�X�#���?|g9��eF��}�����q�^��mh.��3�U��K�?��v{]��dD�m�/�.N{�F���� ��n��T����>�o��>g���5U������C�L��/��s8��f�Dc�Vr��3�����1[A֜��n�#Ƀ���>�s{�_i�o�yld��WE_�=���G��YŪ%�h�o~VK�a{���'!�p��sX�an$�M��q�|>��}�`v�z���HC����#t����Uэ�{�_D�k�Lgu����n�q��z���?<u�+�8�~J��� ��M�W}�x��T�Y̖-�W�$�C��级's�zt5AEO����f��4!^6b:6�\�HS�(��Uv5Fz>mQc~��}�+j�y����C:%����_;�EL/�l(Nt_�X3���[2��(Di�	�%���	���nj�c��Q�kͻ~�y�1��� {����4�'���g�ft�8�&V~XiZg&Gъgq��Ͱ�SN���N"���{��X�m�ׯ7�3�)"6�D�����9&o�ꅺ�!��2�<�΍�@$|�>ͅ������4��~��'o,�E&BZ�'Ǳ��2J�i6���#��>ޢ��b|���ll�{��)�.��>��h6%������Ǌ.�9�.hx3�x<{�^J'or}�j�R��Vr4�}���c�Y	n�#ƭ�36��G�LGD��@��U���2~��ab��j�<���gI�k�ҍpp��}ɹfO���+��D���;ׁ�jb$���.}?�xqխ/B|q8q�q]�u? �곂����[�G-I�x"�OlΞd����R�8 �CA�
�{
d�t�;�ES����1 ���/g��#�|&��̰aǅ�c���f��2�����]�Z}�ݮ�c�AP,PEL{;�h>��[fΩ�l��e�Z����m�I��3��J��� ��->� ~��<uα��S����r�z�7����|b�U��>�����8�]��)��]��[&V{���Cn���tnW����3j$�!b�Dy�ށ��y����^J��p�N_�'9�W_F�AW���t9�ɊҢ�/�i#�Cy���A���ݔa���x�vq�����b���_�G�����vh�A�f��'\�}�[="T]�h��78�Ȝ��H㺛�F�)B�"|��>��y,�M��}py���1��4�����I�[Ej� 8�`r{���s������o��o�/̳m^\ʲ̚l���L�vWd�v��<��1,���kx���\��o��O�뮅*�R�[F��c����ulݩՋP�JҢ�(�ώR�=��wML%,�푁_�.�SHj�M-�!�w��M�q[X:s�Fi-�E]�P����32n)�z�X��Yy��P�:������ђ{L�$��DSF"1�~pK$�݊#���u>ҏrr?o���b�v�*�_�!zd�Ԍ��lU���>'�]%���`}������p�5!DX��������_����"�~�� v��d�md�F�U_�L������'�F`��_��H03�YԻÁWb����R�N����a�$��w�/�&�y�7Q"�.TT��T�	�mjac�>��[ͷ,U�?�s�iy�����@#�)MA���y_B>��w���ѝ&�+������k{��[x�G$��!���uvKy��l|�H�����QÈ'vy�Sz���X�i�s��ck�&;V�iH��^h�˫E�x�÷����J�%��bonP]����/���H��]�ݓ<�}��L��8�_���&�	��!���Y*���x3)�O}u70i9��[�`B��Ox]3��S+1���,,�W���K���'f�'z�N��;�����o�ʜ80jzt�0vط�U����!!��X���^����ş����>�~��,�����w��"B����m���?���2���u��u��4;x���h��+݌�YOc%�;��OSI�x�?}�6�G�2�L/�O�s�>��uu���]�a��n�}pt����P>��K?l�Ai�f�u�bL��2XLۇ�9�9�a��>��c�y��-wʤBN�o�1�0u�c�'�&?���1_H��;�xC"��8ߏ�7h8�'���o���a6o-���Y� �=n���Xk��B��qz��V{ݫ�������;��t�e�T���*B�����?xT��D"����s�s���Xv ��iF�CW-`ֿCҿVnI5H4��յՂ��c"5Y�=�r��|�x�Je��T)�t�T1&�k#vw:���:�s���f�zs{w�/V4u��r���s��Z�a4G��
���S�9\_L�����b�?����C�wg*q�����7�?��ľX�6m��k��S �Dn�(�	��g���J��qI8}�q#�)R��t['�5�Q��m���
"�\�6�r��~�NF��
�-��AL��{꥙� �K�wѧ4q8����"�iC$Ǚ%juY�>)))#����}����qr���@r|�����!���4���r��b��g�3Hag����	�*��ғ�bC�;g^I���GS[�jjjm�{�:�O�+g>�<�H��'��~'C�䭭}��w<W
UHHK����.H:���44Sǡlmm]&E~:�����M�4!wL!�ddg�������$Á� ��~jèU'� �:�G`���	2��O�>9M	�*����2��ax��~��x����M�8kܓP(y����p1m�7"FM��G���.3�����-���ߢ���,Mf�fG4f�rߛĴ�����)���͆�/x>F@@�����\����.,|<[� ����������
%K�(K���<0������ޟj`VωIH���:��7�ӭw��Ѹ/�:G�*���rs��%�ɰ���z�!L�qm}}�z�޸��K˙�D�������KJ�à�sB
�=vQ��J��р�E�3/��Y٣ᘏ���3����r�-�O����Ώ�kϗ��P�(�Lj��υ.F�b����yk���A�k�뙚U���S����b�����[Q�!ZA���G������R�@��3�_�� �1�9�ʓu��Ņ��&�uV�-3�D.��v�́t��(��ֵ?���g��_�4¼H#����w�:Ӎ����rrs���B%t\�Evvv����떑���RH�s�hy�=Nl�����2B���UW�p\䑢�ڵ�����}N���a�^R

	eO��W�]w6������=�p�|/��^�lC�(��B{��U�R������K )*���.kM��l?���XS���A��--d��$T��<V���F�-��bk�=hK|#|>mn�,��v�'�/D��qoo��lR?{j�ܴ*�trrJ;���nց�RhZcO��%l�l��Ĥ�vvx��ȕ ݐ6m}}=��'��-�����'�B"[���O�|d�����3�oǖ����߿�G�|���u;���KIK/���w���͹/��b�e����K�V@�k��8�p����l�7&,8�H�$c
㺂Ȓ n�����|o��]������ajvv��s�/l����|�)<���L��Z6�Mj�h�3R홱%+���G���q�%ڏ�R��<A���~�:\���Z��۷��P��2��VFa�z;Y	пk��>^�:��Y����W�!I^��������GR��'cq4��]OuLLL���<O�@�kM�0��a�aa�|�g�5��ϒ#��h/���D����)S?==��i��~>��ګ����=]�ǝȂ�r8CZG'q�*Vq����G}���A�6z��Ϗ�[`�+Ɉ��7}��������Gs8Y��JI��!Ï�����X�IV�Q��ܴF���لN�YZ�$�-�ʅ]���e����C��I�x��.��UzV"�'�Dn!L��YnO@�����ev&%�8����rR~�����V��ZmE�BT��w��kt��cS\�)����, w������L���G��ۯ��M������>�R�I�����q�>UUq��<�۝.G��c��TB	����B�k��������8[�\}_�rI�2v��뫨`�{��=�pq�}�?xh7+w�����4ɟ�o����������&f`:@^����+|dk:���x�p��wf�8�V$2Z\T��:�����٨�ze��PS����ٴ�������%�tpٿB����۬��
	�^�6�l����3`M�Y����*vq`��˫���g4^�M����1
=�p��I���������cf�@#�g�6�<�O� �O �G���P�p����@B���9�\�e�5��Ԕ8ʵ���.lD[�7�;�N�5w��}Gy H��J�p�@�]@l���(뱶�>MV�!pF����V��?���(	n��)�c2�����͒���o��{|&Y����/�bQ\������	�Qg�h�d� � B���F�ELǾ����y�JE+�N���&Q�WBu������ם����?@(�p'� |�C�oOF�L���j|�av� ��=�#�o(P��4#}oΏȐ��\�t�h����$ )heǞ�!-R�R��HK�'�&�F3�����pO�������~��G�
�PP��'�p����5�z|RD�y�B�2��0��f����H1���������BB���	�q�$��/w��O��O����Q�D�-(�@U2�kkhh��,,�%u�@��'�d��i�2h�|>. +[�5!|,�($Ю���pXЦ�!��!t7�����t������ j:�T�v���%��>I4�Sjd,Ԗͩr}�h�h�35��$��'o3zޖ�T�����&�<)�j�L
ȋ>�΄3yɭ�#-�΍��<��(��$B�����i6Ixm��x��F��D�+�hGA��dX,�c9@�sQ���}i�=.3������*#��>�mؾ�g�O�=$�HȂ2��.�Ӌ���V86B��`�C���}��s<W@� :�V�N�Zm߃�$71���� j�D�8ߝM����WWWcGuI<'�p�f��ύt���/��-�� >��L]hT�2�-/	�^"^���n��Dϩ:u�ҳ�Ca?t�p9=?�O�X	7'�#�����CCMM����Q�vp@�������U� ����geg?z�䉣�5��J�a�@�x 9��LP<>�4� Zr<�Ģ���3�R��1Hq�����q4DDDKy�a�T���ttti�}������			���k�0���&o�ݯ:\T�H}kC�g���ĸ�@�Odh���4���qz�+gF���]���G��:/��2�蕼�y��B�	V�0(˅4���Ẋ��������`df^ٽ�}������jh�e9����*���?�|>*''���yBKg9�!c���(��h�;�c�~�����i[ޯo�E��"##�0�n_.����R�u �q�E8�z���Ȯ�t8������Y�)�����8&I�%<
rӑ��� �Z�}Q��	�ם���_P�b�|�kcVWW� 1����vO�NL �`�oi��;כ��.;�C�
�92���o����,���l}[��+��
��Z�9��N�8�����w8�,p�����{@��W��R)��9���0�Y��CB���G��@�S��,��;½�|fVNę�0�{� �i|+d�����yFF�V,�KɁ���0h6���L��g�?���>v���|$���.���KG��WE����X��Jȧ��		e!�S �%G{�Tp�ȿ��oR9�Uϝ���C^�b��QPdfC���!�:�t��ccc�n��ݙJH]��l(��ՉS��#�Cawޞ?]�A�-q�]t����b�o����.vgK��
O@�[]�t�����IB��)�71�2��Q�lUJjj��Q-�t��(�Y��E]߽ˮ�M�-��&#�q~�O�.+H�0`ٜ��2�P�n`^-7��$;U��ij�b�kA���Uk���X��6�p�h��ugF|�Ξ&&T0R�6B��ǂ���F�/@���߷���b�x�^YY���1]�o�h�`�d�6��(����c���NЁ#�����_��d8��B������S�]�ؔA���Yx�����		]�P��<� �q��L�;���J]�%4���ݠ��+�QP`5�D��D����? 
�������e}�WB�����g�^�ܠ��̞���iU�n�Gm�)� �(�ˤ9���'//��MF��.+�$Ez0�5V�@��灈�
�GIIMU��zC%�+̜��a1gS'�+���i(��?4!�q�� d!�CJ///~�R�����~�����������S��;��������H�l���{tt�ʜ 7������7n'	�舸�$@zi"�_&�N��㣯t����}�\�a<�*#�j�� X6хW���V*U�4� Ã��CNxYXX<_����AaceuHD�M݆b��\O
�����c/[+4/��ϲr���3�� ��|��Ir�j�&HG)0v��s[h�aNNP���s�ǫi�і#��4ff4�M888xxi� :s�Y$JnS$���ÓV��Յ��gi`@
�����	����l����r"d@*�=���@9� Q������H���W\[��l9�~����@>w�G��_456�S���0�ɡ�>���ɁA���٘>���r�&z3���E��`l�C�o��tMV�߇{����O����lQT��"m�vb��k�M��Z1���(��`c^��O�)I��x{{h��L���b^��8�!���򧤤�F�"&���S\__�cEH%%m�
�|l��������s���BE6����Q�޷��� GĊl��5@������9��Ȧ���TⰢ�;cK̍V�oʙ?��K��e�6 ��5�j= eb��kg� E���&��2~*DDH�		�|0t"�А��5џ�M_@��F6�z�����		+i�1:L�<��|--ݠe[�Y����݊����������?ha�Y�V� G���U@9"d@m����D��C�߶�\O�xސ,ǈO�]()�-��G�2�lE[V�gw�T!��/Y��z�{���G��CMO�f��F>�g�� 7H��贮+�Ȅ�8�s9.I([r`D缭փ��s�؏� m���ưe�c8�j ������NO뺡󂬗;���	��́z�['X*""��g�V�7 �ĥ���lT.�?�4{ LPPf���\�CҴnJ!m\\�n�6���ϛ}�[��n��!�15�6k�e�"M�_.~�, ě���+3ib�gL��N�aPN���7#Q23�*2���v'-ɭW����R��ʦ�&�v5��@�q �߂DfZ�7:9�����^���_�ek�f��5C��ԂD%���?Pn�5���I�e����#�b��qR��*��}�ǂ	�8�&�k���LCO�:[�ًJ\�ޡ��������U?�@ A'd�[�;�z[�n�۱�
B^�E��%
��$������ߋ����F���h�&����mu�7�WA���ϟ?S��z���b�V���cu�Y4 6����>m�a(-�ub�E��x\�'&&t+�<!����7�J�[wHቒQ�L ?�W���׵<Ϩ��`�R�$'�z:����B,�ᘵ�':::�Ga�|�������Ǟ��v���ms�5�����~̴�*��5�C�0�􆇃�Ӏܣ����d��S�]�)DIsϕ�^ԉDh�T�r��(==}�����Z��d�8%Q-}�vq�X�B���}��^@l�xğ K@�����BLi}��Cy�֫&��Wkx�b]ƌ1������@���R��w��d���W�64���焄�y:n�'41�}��r@5`��0���eCV�:g5g����ޟXɅ�Tgh8������G82*J6���ƦX�o�@��0_�tk,�q+�.�^Fc"%E愕_,��_���[\�fr,�ꕜE�z���7'����!�E���	q�7���t�48??����d��\�6�Y�	�����UUU�n4�
���񥅕� L���N%$|\�-����T�k[��7ȞQ�����ς��6!p�p_%�in&�$;.N�����MR�i�U�&n��"��N��]��|d�:9��!Z�k������ݻw�"��i��B����w�-� S�?Q���k��k�`E�]Gs�����F��dI@�bb���<���nv��%����n �������v��'��f���?��[�d��+g���:e���E��޾��Y��pp(�)�.>�������e`�Ԙ773���O|����m��W���B�:#>�z%2RR���O�=�l�E$���o����G�Ѥ��:�͎���0�o�Ɵ*I{�:�m�+�_�psts �V�+<k{�c����lk�g���C�L���^�ax���o�		�N\E��߿c0'DF�D�5___�,�� �r��_I;�^�H�����YUU�E�Qb>˯�wY��&����$���f���8�3��K_׾8W�w�v1TpG*��!?.������~>�_�s�Ż?\|���>H_P��{)�9���,,�~����wa�С.�<r��<l	��@� (0 ���1驱����=�hF�|u�]{nb�ɹe�V+�
��Y����6+n���[�pL�y�Jf{k��qXu�N���q�\|�V�<�˗/9�0 ���݄`;��_�� ���r�o���b��K��������b~�vvv ؄�S�[X���� Ϙ�+����o&0�(�Wf� -~��-��Hbr���4�ػ���x��*��d�#o;�a �Bs\ #�j�uk�, �����& �|RrUИ�FzN��0(��, ̍x��T�YQ]f�b��QS��F(��Ҕ7��g-8����0Ã��@3�6fm$9%(r��մ��݉X���֪xF:��`5�+��N��:
����_' ��WPP��{qg�ޅ���B�?��'F�L��Ё����j��X $�P�Ѯ�B�Й�*þ���������頳WKm�܄����O��f��T�#�I���n@�R32�װb
s�^G�����薫3y���i�"�J'�H���O��_�V^OTt�8��b�����o�@Tg�T@⚳@���*�xxe��]��E����%��O��cc��!�N!A� �CU%�?ϴ�%�CǷ�����=1�KMJ0�C�?U�Ry�Y��+�f�%���֏�� H���A�^�ϭ�L&@��̰���m���d�� 9P���C�l��[���ٝ%�S<}*�zM�l̷��ͭ�#k|�����u��_���666��+��fs<W���/��c
�˛��>������d�%��g6�~�~^S��(����@i)�:��vp`'&&��&$#�o̬���z��Q;d2��o+n�o��=��>���I��}�2�g�**ßk��#�������ʏ����ӧ���]��؈P�-]r�`�L�O �P�ũ;�_��2��������}H��N�%����(S ��{���~
���A��ҲhN�ҌA�L�|���8���hy��S0Y�Z��`o_�[dH,��q�YW��uE�����&����>/n%]����jf�&���x}������:.�f��oѿ����R�ZG}�3K�ү�4�'������ܩ�0� ���z_8��+���U��x���˴y���`o�u�O�b�&Z�Ķ·�W0ld*�q�zT����x�k�b�{P����j����8�j�!P|��q�=TXf���rA��*��p�i����g4�Z9gK����&Wi��`���&4�H�g�F�/�k@�m�	~B%�4bb=1�?��B~�i��m�]5|����\}�* �ibz,Z*b����E����뇱����憆��M�bI�Q���C.%7	�^"�q�����ђ|�g�]�P+�oS���������IO���L��3�����)�JF���U����#/G�xI���\L-���䎮�i7O�jFH�0�#8��PᆞO���Ѧ�;�R����_Fk�rW�=����E ��D��h0�t���ý������7�E��<�_��:	��t-F�>7C�m�Z��jA�;���R�L�cT�����w64ד �6ѭPԘT���988c*^^m�B(�ʓ�#M��"s�Q�:�ڃ�m+�n��ł��k���ݔ��A�y���e&!%�S?0��WX�R_�il�TK��Z�+��[K���}Hpٕ�|�]�ϯ�]����"כ�u�;�bl�N�oZŇ �ߐ�|%2���1t�]NMO�GB'��*12�2���s��o��l��A��ښ� Ӑ������������rK����Q��Q �1�aaaL�D}��S�憶q?&!����=AF �=m-�D��F	���ԗ���{g3��%��%����LF�n���.���Hww*62���nO20"~ �On|j߸���L�w=����aS�"/�r�bhH����q���x�� �w�IGy�ߣg��C�T��
��l�X��H�:�ez[I�x'�aG�I�j�L�Ӹ�𨩥�^��$ccc�ü�J�<�[t�Q��po1_f�`_�Nට���r��t�M",K@$��⫻���3j��><�z�x��d�����S����ם�i��KRT��'���[Zm�ya�0/������u��;y����i����
����~W�89���&80�drddda�B=*�5��l���_��a���s���˦���W
X�q�PV.�V��͸q#B�Q�k�� ����KjiM$��4�9����1t����INJz_m3v�8�D����7��\ۅ[��Y�GI �}������W���I1m�����q/fǚ�0���2-�ttL6���+��f ��֚��ob}3�����BB��;aX� �j2g=��B�҄��8\BB#fQ�HҎ{Zl2#������`����{࣑"#�X����`����~�Xb���!M�"���A�ؗ��::j�lTT��^0XPO��P�2�����~�_��A"���z{����.\�&ȯ���q�5E+�ӷJ&���@ǫ���]#ޛ!��ƅ3��z<����t_��:��О�\`�������S�E:���2�'�xx���{}=�w�:/9�@�y���+�,�0_kX��ɉwp*m�����36%����A
*��ȣ$Ez���K�򞌨����0�/͵���Fq}�_��,�[@Dt�^T�x?69��\�du*�!UR-b����x��e�ӕ�wvԌ����Q�O����o�)�"�H�X\R��%P���6wJ[>��dMD�;ЏGӘN���-9��} i�}곐���h7FD,��ǣ��?�(b�b�w���f�oiL��l�e��������9�����!t�S��*�')0�0 8����i� �c9�O��n�F�C��tk\Կ�bv�t��r�U�����9�n���ng�>Y����\�������@� x��$ޯ������Lc #��2�Hgb�h����X6�����@�	z��ό����nw�!vI��9�)k=�_����-��-�(�&o��+��4yrA�=O�^M`R���!��u�2�.�x�yJ�o�m�s���@���<��6P�@�����kf/�#��ߣ�4�9�D���+�^z��ѥ��� v˕%%%
}?t�;K�N��3�s s�O;�] $.|m��Qu�UPZ:lc#&�u�;�H���k?�$
��cԴ��#�m����=��W@� ��U,�sx�\����2;{D��Ä�Ö> �)�1���`��UgN �f�R��x{���~�M��޹��r��ʅT;g^u��n�N`$Tq]�n�/���[d}��i,�d��=5���1�qVTy|�T���_��y]�Z��}x���Y1��y���W��a(1�U���l�rpR��K��X�vp�)������m��1�'~�c�񤦯��-�F�C�Q�ٙ��@2B�8\�.F�r8ȫN� G��#�$��M�K<����=��rM�ߤ�9A����"�k<b�F�5���.)ybhh�{PT�3S��) ���v���9dvbC�-��F|���s2�k/͝�S�j�ÎD��ᦱ<�UB�:��h9�a��j<Y��x:�������)oh��|�Uggg�MB�k-�(ٕ���@`�.�r��|}}w��/dЪ��+�Ѵ��[{'�Q9cK.��o��uvVVk)�����7�B�ȈT��t����i�B�33���?���Bb�7�j�s�=XЎW��H�ha͒h,�?P���ֲ�6�24�C�)�ޑ����&���L�����M�Ƒ���5�W^��U���}Y`�S2t�LYw2�ё����R2�v�`g{����_�>>��Wth�����e�T�w�Bi��h��Vǧ�|�y��B�*g0���J�їn��h2w%sYfM����!}a}TP@�4�Xc�34=3����*8:=�;�nN����	�u��4��K�Ĵy��{PFJJ�ׯ���V���&6���
gS����r���[�j�`���pO��.�S,7Bs���!�[�%X��~�P��J�I�,��n��/ii��,�<��y}{zĺ���P}�r@
�������)���w��Z����������[
��םKGO���vi�_�h��j�<�l
��t�� O�9�I
��f�1,\�%�2!t�j�{.�U5){a`@_�~E��",z���������𘳯�Y �G]���0S�R�J�1*�o]��ݩ4/�%���[��q`C�8�T�2X#}${��t �c��?��pssgegSQ�����B	2+�x�jV]�c,r�����ݯ7�f5��ѻ;�"ޖ��
ӫ��_2��z����ƭ^�KC�y�%�"�6��ǩ����s����z0z_��P�8F���tL/�D�S��|��MUC#�")#��R�%�|�]�H//���Y���7��$�]tkl����������qm�t+��h�SD�����%�uvu)]�K:;;C9��qޞT�9�\�B�����_�|��!x~'���G#������Z^~���M���,(���|�
�b]�P�׹�H�[xd`�#R1��\^�k�]�+���UQ��+�xK'G�n`�����⪁��]�԰�;r�#%%%9D[4��Ԑ���&��֒ ��Z�76���+�3Vl�vq�JXubZ��� ����5H�����Κ��H�	��l��3�Q��*)EO��:�-,(󠠠���Hdr�a���c�-����#��� ���Uv�9:r0>�+..���MJ�����+��ׯ���FG��|E����JF��$LM����E�jkkW���Ӻy�g�ܠ��<�ƪ���7��q\�DXbѝ�ﶹ �[[�_��dt��E&��/��͠��e� �&y�rѾ���"f�?q�7�&M���8�#uP�n� �E&=�5A$��j
7Y�����V
<���?0���sZ�%�?}�t����_�����C��54m�9!!��:�;s��4AT�ә�Ξ�ܦ�9k�l�pF��x������������ظ�A�(T���-�Z;b�ޟ?�PPE@��� �� t~-�B�:�s�]�b|�.6�OJ	����2��Zw���u��"�B�㵗-��xB�k(y�L999�����ά����0`o���G&��ΏKK�HVDNVkk�8==�:��?Em/Q�e>���rG�H��$m�y�_�9�]��r|����s��ҷ���ͽ=i'��443'�q(333P%��:3��~.�b����7
��������	��|�}�N��`:������<@ڞ9�Xl\]��,@
$��~l��J�uY��NAދ���j���6��A2n��s6���b��[��{�\+��gl3���TU��f���E�'&�l�TTd���:�^�$�Sz���_������>J{0h\�� 3O�XĊ�n��]7����(�P�O������J4!��x�t
_L��Tk0�(s\�A_�q��/&z�I	Q�z1f*Zn_0�>��(ς��å���}�};����e9��'�G _��6X�swu-C\���f���;�pw�;<6���+ُ�Gu�SS=�m��E�I����D���"#ш��C,AN�A���;�y�#�ƞ2�~�|�~�T��r�!��>�EÒMʎTгD���\�����NrI��^II!v���2�[q��t1ODno�pC�����4V�E,_����i�'&B�9�ҕI]Q�����4�͛V�4��N��F94_!��A�
��y���:�	�iv��iZ-���̺Р#=���Y-��`�b;�LI7X�K��_���C.����(U��VQY��3(BO�m��8j���K�:v}���e,���1����ՠ(��&J-�����iY.}&���r�Q"�W6������[��f����_IC��{��=���w�W��-f�����=����K��n�����{���?C����	:��ɩ\G��Mu�:R1??t��E���g�z��3�\H1ç���/��Nl�4!�p�����dօ��
�&�[ ݵ��O~x�B��<���x���N�Z��u� ���Ԩ0 D```�.;�A�M���E�^U�����I��^;/l�P��pSdK�a�L=TF�J�	?���tpx��8��	��;Q[�������Q�\�M�O޵���PS�s_��yM-1�z6RQ�(B��>lQ��S��=1�/x�a��� Gˏ��̡)ޟ^�Fn�h�CW�Ʒ���z�>Z��E�i�ǻc8�2�a�'�bVi)���^�U��	pG�´�_���[�!�/3!X����::���N�KV4'(�HV�ZR"� P�`�Adt$:-.!a�ɦ.�m�$tB�i2t��\%H7���>�ؼ�?�QA'Ï���~�Ĺ/:0�>+[��-f�CT� �pZ9Czxo�9��v٣�˧65�/��'D���k����dG�p���Y�~�I<�
D��t��!ظ���e�[� �С����
�d���L�y=P�)������tYe�X��EA,M���������k���׊f��#�����#cc��琍e%���9��������k�n���F.! ��-%]�!p�)i���"��H�tK}s����u��sf�<1�g�I�����p5:U㖼��^��(��_�~�UM�]`���"�355���dė/*]�� ���O��aY^�]y5PYZ��hv���r�{-�O�N��襎����C��*ދ���
��,��K;����-Ye�����/G����r���鍓��zAJC#�f�J��
�;g�I��Ն��h˟���9��C*L���YB���kP@P�}�f8᧙��b�0RM��u����ʗ'@#��9(**���o	�WTp&�l�����}s�t�2VP�W�?k��yK��0��;�ؖ�ZQt���/�Wz�@,�r�}�B�_pIIQC�	wqE�eU��rφ�[�<<=C�ɡ�L�h�yн칳3O�{"BX�TH��Fz��P�D���
���_�`�7X���_��~�K�8�4MMI���X���U�H��4`?�8\!��	��(+�����51�����"1	I�:FI�<����l�>�� )�N6�.�\� �u�������ɫ��W��2��ߊ����P�W,��󱘚�w2z=�u�<��*�P�z51����B��{ ��9JN���ʺ�����5�e�d1���Z7n�UXK�� �!?�67�y	�f)T���	�2f+77u��>��Qr�>�P�` �{xE��4ld#��6�����z�����t{&�շ<�8k��R�͞����9`�ґ��'�b��`�� ?�-Y�s��U��,�o8�΋$@ђ�$���� �P���+���=�Bn4�V#��xef���l���F�Y�Ğ?y��JJ
*E��/�_��yd�J>(��%t����/���\�:Ɏ����1���H����� $�eq-��>H����r0+WX�����g���iY�)�d�eaa�O@���kH!�������n���f'(���� 'J�5�aT,
�UK+0�����Ӕ�j=�iZ��������BR����ٶ�m�i��S$��1*F̴E�@��=K��Ҳ]�EK��&�ҏ�kzc\a��;5��f��74ނaC`����Xn���zd>�?�T��H�"}->D-u�N�ʊIL\\�>��+����݌E`ވd�,,1����*u�7��.8?�@�Vt���e����^�.Yt��Ȝսi�%�H.b9�����.�?�DlllCccg��O�<	G�RaUK��X1茈���A}X�����p����}��*���O�G,;�Yh�'�m��Q�X2?�Z�V	Z�G�p�����\���E%�̌��<�߾��&����D� ��!Ζ�#�k� �@�8��Fj��%k5f �~.��� \�/������]Ͼ]O��*>�3Ʒ����k��OX����s�r�Lْe��ѣ��׶X��_^�Gٞ��&��G�>��:M.,���(�9w���	�!���a@��?0�o\�Ps�Yc���gt�.x{�����م�P����~8����@7��i�rdl,\�����6?�/��2@5�tuukz�o�m�=��a�cm�/eś���B:eA�BZ4333��-YI�~dÍ��!��L�;&..X�Y��P|)5��2$�I	@�
3tI�Ym�	k-`z��|��H^�E�}ySPR�=��d��������c����������c!h��b���'�B_T��䃝UE��+�R��z�|�ӝ���>%����7v^)nݷ�C{(�s��������dzI!��pIV<϶рӸ���ܝ��{ӭU�@Z��"N�h�f���I��$}�65uW�ʺ^��D��qM1�-�7o��v �'���阮�a��N{c���;�e�)c��w�(@�̼4�us�+�ܳ�I� 226nP	�#n�/�����V��Zss�O�Φp�a�z�4@�B2�Cr�n=�����jo�d�)V����0
��)*--,,��ZJDn$eif���ðw��RNE744��x_B{Ҩ|�����e����E[g秆���h�����P?�b>���J��(hS���<����Pa�$�IzI��D�}��������_�p�A z�''MiH�8sDD���0(�??�^NN�Q,>��uE=r�}??q���a���j��E��x���� &�p��&�ɛ�����[�B`񹸸� }��_#'v��ÇQ--"@-M�Q�}o�'�6rW^�W�P���n�/����^�n�w��`��9w�ųVk#�eÜ���+#
+W���W��Ϸa���o4�5���M�)A�:��gC.6W�KV���8�[H$Nk��\�.�K�Tj*r�Z��5�-*t�:���޸̂�$k���C] �5444#�t����_i!:�`+})%��i�Z�Z��T!x�VSx����f�V�����S_�0�[ܦ�:�??9ʨ������oMM�ݪ	�P|z�������8g��e砱����M�������q�K�}�Ny,��� �U)Ӟ�<���S�S��Q"æ��S��m�����r3��e��p趉�:B�&G�F�8���B��ErT9��{��4�U>��f���ݻw��$�kiK���,�ǒ���0����?;2՞2'�/u ����܆��h@�-�If�sf��U𥹹�����	 �x�F�s7����#�!aT�T	�k��PXK��&_�݂�K��k0Y�N�����0}R?P�)A��/E����^��W���	[Ђ��S�F�gŭ�QC�֖{�O��ô���;`a����͕-���蠖i����w�-)i��f�I����OB�ٍ:쩐���o٪62;��J�c���2�"驩�J����tttP��!��~�'A�et�g����Nq�6�|Lm]�<ݯ����J�rϹz�i�Ώ1���M��M|}*���S�"I�iד��ErЕDx`����S��� b�MO3p�Gs˺�����v�N<>xF/@�z�����
�+�#����x�&�_�=�E)�[����g,�sr0��ӆ-��$�x�6=}��D������W�bB��X�Cjhn�z�&S��R̃us]�0�������Q~� ��t��ϐ%tBt<E�;�tJQ7���4�$���������g쩚!���V9���.nn�Ϝ�`t�M)��d"��Ɯ�}�]�\��ED~����@7��>�p�\��E�����<Sr~A����e Ƥ�G�������홀��3����y`t�]u��K��S�r~�����rl؇���Ұ�WT4�V�]�^�$� �|��&<�X����l�Je�ς�=�ۂ��2^b9��e�EpGFFj�8�ْ`MdQru+gf�o7m�����%]�]��fZ�N�`c�hDF��7�c�U�0��L��_�=�z�;��v55��P�XS��+ί���Y�^�MHX�5���y�~���o�B����&��+�xZ=��)�>�T�� ��r��[�PgG�tt��o	˗�Ap��Ąe�du�^�}�{��x��T�
NN[����ksH��a���D�{=ލ����i[�p��A��'n�*V�vg5|�[���E`�L(�6Ws��}�76�U���wu�^�ZMfU/���u�_�9���������؍ F����tt-�Pĭ�h������
�"D՚���6x�3�o~�c����j�[c H�yXN�H���
��X���T�~���Q N���S�.���-� /v��F8�_Z��9���W��^�E��
?~����IӉ���|�̔�{$��.@�M�P:xi]�F���m`�>t�I��iE�.@��r.3�����/ے"Y��
��Wj

���n���&�1�î�s�e3Tpwxu�����WH���ʳ����/)))T�'-^�����dT��ײ��̛�kkj��[u�חp������~�AWOw��S����ZK�H�V<�c�jaq:6�����`V�%����fx\�|l�I���M�P��X�܄{1!���6�L�;9��"<wdn�x<S�C�v|�ܹ��,�j9Y���}1�>@���Еh��q�_����V��OL뇡��O>�7h��R�\����js�8�*�2�@�=
���@�_�!�YC��~.��Q!:k@l���+d���9	�/���UtBa�v�P̚�O� Q ��-X����qf�`�Ϗ�>�^>��ppšvd�Ǳ�����i�*�uI-`C����~���z����U �I�������Qa���{���W/�ii�8�A<�x��܁�P4����0X0��N�pǔ��攈(;�Ό�/Cg3��\�cQ���ڽOEN�	�j�ӟ�
���2ģ޻�u5-�~*�,LϜJvJܾ�O�#��e*k�
gft>Lg򫪨D��&��'��C ��d_V]�`@.��DCr�+������A}�M��l��������n*܈���7K	���~gz��Q E��prZl�(�������Hٙ����}P<�$Y����a�)疠�����-�k
�]�f*m_�Zq&��q�Ȼs{GxB����Ůg�[�w�BuV�@�)} q����'�
5N�ϡ������&���kZ���FzhN���i;�{��3�i�����h%[>�bH2���;z����h
�+�T�z�%�������#���I_b-���b�qG����o���,��N��TT�|t,~ݢz����;��Ö|�;�G�{�ZZ�����h�x���P��9uC���;�� ��fz���>�H������!V�p��<*��N͜CFvv��c��ķo)�-��_����}���Cu��y�ٙ�$���� �� �%�'��Z����>���]��ô���������缽��k&�ϊ̲:n�[!ʻ@�:��')���sp4³ֺ�;��{��X���uV�����l�Z�۳������A������*�x9b��=�YS�6���C����#�mƩp����_��?9I��N�0q�\=��@R
�/����z���t�Qs@Wn,:���1�<#��0}�������m�e2�����څ���\��9�z��4����7��A9Kfn��Br�ۅN6�;�Vcx
>~����:��=��S�P71�==PK���8j���e��KIF���LY�7�����p�ќ��x���i��ΞZ���ȠR�N��Q���F�t��L���j���Xx{�(j,�<h�����x*��F�9j���uL����J��k�x���#�l5�P��z�&��$���N��y�������e]�Q�X��ۇ��e�:�)��=o�D
]�r�s�˴1�= �$0���w��&�ޣ1�.�5��ۯ#<��5E��?6�˜��vu%P-�W$ؘ���L�|uy9�P�sR���#�1f�� �J�!��}�A��פ�:��Z�>����
8
�a��O��������<���V-]۟�}�VRR"�(Y�bY�\�b�����d�R�Z�<vg姙0�(JOK��a�]���~[\��z���з=��q�n!:9o�8���ׯh��D�M�8-�Z�?|x3���:*d���-�8�k���O�	��^��D�Cw�y��aY�4�WW���$+W��e%f�����Ee��ͺ������n�x������v9z��/���.#��׿��ĕ|L:~�㺏١KI�h,�IM�~�����mc���]3Kn�o�β���|y?Wy��f�,(������j-�e?`�jJ��r<����wa$���*s�`zg��TGECs�80���Q�=R*R��K)�ki�;z�o�M�/�Ԗ,NBB��GYB�������uW."�ڦr쩫+}J��kJ��ѣɥ���1B��3\�,���	ئ�G�@%� �{ޝ�t|ǘ>rxZ$Y�R��i>,R$���ߔrU\��F�1���i;����l����!��^�F��#�����#��h �����P\��a��ݳ�D'ѱ >0�VKKJ���<_��4\��N/V���wťǂ	�:Ⱦ��I�&q��u������σ�����|�fv'5t����� �RRO�������4>膳נ.�Vij�O��t5�z3��УR'�0C��yfjj����vK>};����M��Ö���C�Ԁ�KJ�:|��	`G,��N��9���;�R�u�-���y�M�_]2�v���S��Ӈ���(�<�f�T�b��J���?��H��D���Z�H��"��{�^'���fh��8�t?�����3���/�	Xd�t�_��B��۾���A��dKAh�D��&j`hXtH)�����PCW�猋�55o�qE��S�Vg%&��P�yC��]�����~����Jn`� �x��X̬�3ml|�A��DS5l��-L���o�7�}��' ����i�Lf��utҎ=c�X98�E�W^|�i).f
|0�����^��*��kER�|z���� t�/z�"n�l������?�0�΅�r���i�(���;\E���Ŏ�#�l���M�l���#��·+4 �]DR��>_�:f��[��
�Y�"q��ޝnHxV�7��&��a�z�=sC�~�{c�)"?�8��<���v����q{'�p�� DDD��V�
���N*...��<v�ɹ9�j ���=�5zV�OZ_r�:Z�&*Z.ޛ��5�yțf������ �I8���x<<r�$PD�c��]����]�����3��o'(���TT���w/�uK�+�[h*su�ć�&K�(��0���|0{C��i�E���8T���������tS}�:�ď��3�*��q=<<�F�v`�)$/�=G1ɘJ��{��8l�l0W�6�{���~������&�(��ҙW���z�� QNq�ш��Z��U�}��$�����E�˪u�Td�}������.i��q���������3����_��'c��$y�#�Ҟ����ͤ:b�b�j��P�� �_��;|���#�����6D�鯬�K�D���O���L��]�M�F���Y�������CA?�̴ײ����KN�!����hV�?$�z��FUpXu��! ���$E�e�}� 	A&�W�[6��(�!I:�i�sb�w��_p}2��@u잙����� 2¿J)��k;m��\�~-U#s<�'�_�����3��	:����������r�W����l��~9?+�j���(d��X?�]�(�S�o΋-�(/L�J#�Pa�s抑l(mEǋ]�w^3}@��J�G�}L�O;�Ah -Qi؜t�
�t%f�r1a�z���KhUa��C���:ւj���&ў�!��6:]�??����:昡c5���T�h��9	��.�'+L�x(nh��Ҝ�E�:�o)	���ekʒ�l$$� p���R����������pc��E��w-D�k1⎍�E�ʁ���[�w��}�,�3�eX��A������Q'�2&�&���iw�Q�@
|g�K[[�I���Tz�Z>>cbbؖ��gz���I�;�����òÝ��ɬ,Yb�5�T��6�'�#�r��o���b�mf��AԖ�܌�|bq1 ח�1���ܴ�G���[:����(Q�+�{;�Q׉��Rl�B�߾}cl̰ G%�y �v�ݐE'���B[gԤZ(����5UY��B�=p�'i�
���M�xf^���߯�E�h��9>F��ϟ���٪,i���c�-׺�nx�M/qN�Hn/:��X��MJ?_�%�o��͂.M���X^ ��K608�va�v$����>�>K��#�4,,,Q2:�;h�qpp�����Ġ��d���~%��+Q�"����h������IH��c����Z�H �d׈��^��A�,��Z����s=V��O��4#u���w1V�������/#ؔ���o+f��e
'ѩ(�|�44���33�A$x�<��Z*���˩�b��I��3a�S3��G�|Y6��y�V��2�e�y#j��VA;�݉���Z����o�E3��]]��{����C���KC$�t�v�AD)x�Z���łQԫ�Qdl>��j	?���J��0I�9=���L`�\�"��ȴ�H�/lЕ��sLI�%���/�2c��-�Ik�8��ٓ��^�b۵�/�DAf�/UC�����Ęϗ�m]��)�����ry�{6@�A7*]��@}ɑ_���z�4R�bn�����^f��ѡ��|i�L[��i�;^�xArr���~��V�~�v�9�?������uJ�bؐ��T�ޞ���k}�K5#��쮇iv7�Q�٠z�������%V�UA�D�듻%EE�zzzB��q#.�g�83U�Ա�_SZ^E�V���Sp�����?1�>uÝ�� ������V��}@i+�D�q���c]�qz}�sܞ��Z�mS��%�w��D�l��.d~gbgo)5���k�b؇8������-a����,Clu�D('�{V*���,�j��x�j)��!��ϵ��aЭ�`�F �r7�pC����������?F~ʀ��V�g�'u���?Y�qkw7L�|`y��<kM�ڕx�=$����q
"9c��S�ښ�O�,���2ZZD!=f?�IJ�n�����'�c ���3�������eK�	>��b�4������kE�:ߏ�sP����$�������Ch%u�V{�W����Bf~��l4�{��]�C�!B	,�#�4�NJ/����1��u,�W�?
��L��޿x<���gL`�����i)G�V�\]QA�/Q'f5��w�A^ �9��RW ��^�j�#�U�D�V�ׂ5��C�y0�D��{��4������Ъ�=��i�p�V��g���fٓ!~Iɜ�[�a^�P& ����R'JT�t������%B��;�'a�!��j��[��.��Z��~��s�\�r͗�."!ݷ;��frQ]Ŧu���iI�PBe���\�ɟ��,|��x�)PѤ��ĽaXd'�R���W���LL~&�m��v#��+avЈN.#@!F��ٝ���P�ڜ��Q�	 �I ����V1�QcY=�,�s��|��	s�{�%D||�����A�~aGGG	w{^�Oh�?E�!x�}}��9���0ɟו���kO}y!�&�� �&+{�}E6��|}-�ks���3V�;�\Ê�v �����[gth̈́�444��;�Q���nRM�qķ�������UAr�Ohy���ѷ���w�>{3`�!u���ݹY[�:]�$����a�Zr�u�y�D�w=N�?s�,ہճ�� �6q�YA��i��{m���Ǐ���,�8�3�w�$����\�j���,+Ø�%����T2Я}�B��#������GL�\�V�r��2��x��g��@���5�녲,K�Ŭl«������BYRHːebggo�����jd�pJ�۷��>���_aa�K�T�e���[O������� ��},����*\ =.�Ѕ�}��I3�M����s&�X�Ԕ��D���x��.�[���ѥk�\�=Q`;x�C��.K߮IG�p�!��R�D�k��� ��\Rg�����|UZy��zrr��P�Ls�+	�	!o�H�[�3������&�)0��E���OOO�g��{�N�����!W{�xH�RE��bb�Y�9Z�Iq#\�Մ2K�d˴C�D�fX�%jo�L�������8�\�d eB��,���	;-(����]={�EI�w;���#a'��l kR2��,�Sc���RBqi��t E�8/u�4���umy��������|۽�vR�'�y����t�''���;� bdk�˫���-b�i�{�Xf�+(�/����92�
n�z���Ag��BEEu�5��*z����1vh���ы�h����>7IkI0��@�,�|�j���-���A��T�YS��Ю\5h�����V���qj6�(�v�Yc�@AII8�H^��u�Է���!x�*Ic%;d�ux���������?�p�*�ɽ���5Y*�P�c����߯��r@T�I !-'�n%�b�Yki@477Cg%�ޤ�� TkeuM���2B��v�tv�$k%�9X���[�B!{��"���G<�㸷�b�x啹�x��8?����LKKk�=G�5��'�a�2��.���_ٹdQrЖfYY��q�SrS?𬭭��ۼ���. ��P"���0:�[t��Q_����j�WHH���.�?4��777Ho����>�z����F<��'�yL��}й����й+*K��ǩQ#х�l` V�=]����w�����


�RR���+T��@+$�~mus����/���P��*Z�(�6�����F�I����!+�@�����w3�e٠ە��?g�[���J�s}����u���-k�8(�@
��R���>�8;�lhj��^}^8	e9�ۨ�?6�4��G��Q��+4�J����s�����yE�=''��^�R���q�M���$���e����֧z3��''E������~��*[{{&^Q����DL[�.�o��7%���+�����<��6ߌg�둴��!+J�u%�kbD��[����	WdLRm)/�*���$=Z�	�[�h#-�du�Q��.�N�jD�q{��>:T7��[�A<{&{��;�AĤ���J:���qfmc�OEg�?�s�*g������DF5έ��ʨ�9(�E=�⥺�5��������1����]9ey߿߫�^̃`�&Ib��b<W�߭��\��g����vj~d3���=����l� ���]Y0�׀�^�0`�S ���y�[t,���3|0�����MܵD�n:�����-�2].Vb�|i�?��3�DZP�cŗi�! �q�Chs��f_&��\�Vg������d�V#Hpux�*N������;��xr�/K��Frgg付��Eȝ}��B]��6;���8?56�ጡs�h.��;AG��p�6"�b�N��y�"#��ͫ��޹\ʑ�/h�\����=�;��Ry<���;;b�*+���d����v�k8c��.5/��r�za��*��4��,��w>\mmH0��k~D?��<������ qy��>=���M��$�����w4����צ�h9�뮿~�d���@��BU-��Y�1WVbZ���g$�,�z,j�0T�������A����"B�ⱝ4�O ��gۄ�ȱ-|}�v�`�l̫��e���B�˰uߞV_��Q"�$�S�Z���0��-�_���C'��*>|xZ7�'� &�K,��N��s��z�kZG6z��K��!��.�>���n��!� �X*�D�GF��^���1�C�s����b_��5�c�&b�����Ku���i(���_.�'^�W_�-�8(H����=:�3�Wк�h0��U�ѻ�v��hit˺y�>v��! ��4�Ö��m�`n$��D���B���bƭnLo��q��߷��.��� 7�t/��%��*�h�`�kI�I���gj��H����*u�LsWM�P/�w��	�5׺�Y��5��XZ޼4�#�qbRa�:Z�;=�j�h�]�7���K�J�=�}�L=�G�r�ٔ�:�L����kj���#3^؉���iD�
)�Y85��M��
��yt��]	�u��˂9�n�پ��A� �S��2�:s}̄*'���D)��ۃ��y��*վ7Z�8���Y�gT/�Q�Sp0�6ġ=�����||�_X\��/�����i��X�L�`o�����K�5�~x�
����R��3���ggq�A��A�WTT|���n#E���$��M��>{=�w�9a�ZJ$����V���l5Λӳ� �ۭ쩘qqq�ʠ���4MN�t�R�<�|2ߘN�]M�9���v�_��mβ��EƐ��̢�y;�8���K %��W���M�y��t=��!bQ�uӡ���eE ����F�{Q	�����\?��ϡ�+]��c�ݏ�S��@��C��K; �����]��E �[�r%���3;N��Db��-����lM�c?������uVn�����,.~ہ/�z�K�ȃүlm�o�V����?�@����;�2%�]�7����P�����:{��G�xF�-����3�e���X	��+� ex�̧6R�UA����ļ�K�<ENLF�6A_j��Ŀ{G�Ņ�z6fnN�eq/��Q?�}����J/�	Yt䝳�f=��-Α����^�����B�w��%�����E�q.�(��;�]��,�e��>y�g �*���:4�`8�,jh>+�ߝ����ڑ��zi�*�Z�w�/+}p#^.�<�DcNT���sMTD�N�⚌�+� <q�k,(..��5�Aŧǝ�6Et\�q��=�o���cyV�:59=-�������=m-��/�kh�.R�d�
�^�ӎ�$�|�%Fꂖc_�Ȇ�R��~�������E'�i~Z8#d�<����xUۂ�y:O4u6/f��R�k�阘ɱ��3�32>=���q��0��f�釪�_���,��7������Ap4W754��`Z��v]>�G�#7�c�:�+��z�'J��rߊ�u��P'^������`����֦913�Q�G��c"���:�/E���%�gH��\�ұ���r��ʡ����ޞ�B+g?ά`8�ȱQ�L��g���icƯ�G�ᣣ,z�5ϛ7��k9q��>�����4<�𿫨����� 3����-�z��e�dnK57�r����p��M�[`��<��Qb��m�ʆE���@	��Ę=+.W_ Q���iR?H�L��[��N����-�`�!Sġ�w�=FNM=���O{z��߻On�:���||7�nM3��0��]RIH�8[�OD��%''����MX֚�Zg���i_(X���%�IE�!��"��@'J�]�cQ��1����+�'��Ȗ8��C63�% ���&X�࣡��`�J��1���i:���j`��Yֿ��n^���$��c��U�;#����㬞hX�r1F�j�=�Չ�����=��#���Kd%_��&���:��#���3g�70t{�c�=����9����L�_�ˇ�Oi�F�\��]�/���	{j_z�p�&y�T�������}��1�P�{)�����ԁ0��|��i��)�Ğ>�s�uo��m~�(�'eﲲ���3�Kb�A鹶�@�X�ɔO[E�]n����]?���PP�������/�~Z;4��D����������E��H[w:���Y{�|(>�(�JR0�z��Oh��ϯVίb(���Wl�<6��z `a�6%�8U��������Ķ�6��BB�ѫa�]ɸ���bZ\��'�Z:1��+]�g�#uM���gwHF1�aC�'
'Y��(��toe�Z��Ó�؞|��
�4�c�\�ʩ5w���@���m�A���?��T�\cP����v�\��Տu	r�����qc�ٴ9�'C�)�e��E�/��_����7ŗzl��3�g���/7ғ���¾�r{��3�������c���*.X��B����%� �Нk�����Cg�u�`�ն�(֯�����-�䖺��n���&H���S0�8��u�{q+���-������A���{��"}wL/�����Н�!m����s�j����.��5Bk؀NJ"�3�����/)S��\qk]vk�ih`�>����q9�3����_��t�Чubb���P^������I*����!h�b�����W�ʖ1���𠢢jq�P����n�V����!;�Ll�u1¤�F� w_X$*�}bŠ���E�걑nX@���(u57+��������>K��:h�2����,��'���V�Z�265��:�˴ш;<���s�&�j"K���K��aa��5�u��BW�6;x�*u��u�b�����޿]!�	�\��ɿ�)��)_9��}�i7�*�z��^���GLӋ^2LJ�C���*	RR�&&u0
�QM�c	N�Ύ��$���ń��O���|�UY��f>Y�".<�K�[���8��	�47d�Vs"'nW�W��,	ί�/���ȴu�������i
��ؘ����2-�����
9{{{��gVvv���?TW/�.8	W�t�C|Pd�i�8�����FA
��1{h�5?�*<�������\�x$���sw���b�Jsp,۾i;��Ǻg�H:P�[��Φ+eDk݁����~@��g5���lX�0Nt�诊������7=�5�ž_8���>��Gmn��7��cv���P�/�L��P�.w �9/L��i��.���^��p�ڇ�ʰi;�"o`��bܤ1=��}N�/==u��1�`zzz�z{����I7p1m-������@��Ǒ���1��i��Ɔ��/9p-�����e;y>�B˺�1�a�����ۍ���.//�W?�M`i�Q�����[I�TgO}�\�Ph�O��髟��=��E�{8���D�ߙ����X��p�O�hk�����O��;D<-��h��Q(l� NP�������E?`Y��G����B����8k�8�������V�^566*�?�;�z���o�}������� E�.h]�i�h����..5��|;��p)���GG��L˴���7�'c����n�ki%��O.ӭ*��rB���b�����U�����9�y�$�q+q�?��:��j�iV�����V
^����|F�G�)0�RKdL�B>�<<��r I��_=u��e%�<? �x���!���4^w!�'2|���hu�|��jƗy1wbƋ��П��V�BY\���|�J\�;	�ڽ�����q�?(ʒ�.�k�G�L��ǕŚ@J�A{��]N�6v�K��=R�;.[΢�K)����a %ب�M_�U|��ӿʑ�1ѯz���������{�ߎ� P�}d$� *����9/�� p����.����䌅��v�E�N��p���Y� 8�Ԍ�(($D��D�Zz��i�z)/� �F��R�Ƕf�=&�^�] 6��DQr�1!��pv�,�Q�r���T�8'A;·���<�@����t��ÖQ4�S�¦��l�#`�.6�BT��|7-G���?��j:���2 0���$��f�i�5ٰQ���g�p�<��~�Z"^J�X;�F�@!��HC�Ό�[�ߧSnfO}%�NXƼU�qJP/�>��vcr�VpN%L���������$�$*2n��'>�WR�)S���I��G�q���߄�Rq��aX��9T�?� E�c�ﾻ*u38$���%U��ܮH���ݓ6��B�{�1�Y�k�5Y��n��!pS�Kx��% �w/��A'��\�:7�ї��҉/*��T"d�h���מ�SSI5x� V5�1�ZGZG��2*Q� �8G�^L��n��z*��M�0GB�kߗ�*u�I���Ǉ�@������\�9/ܨ���Co���2�	�0{����&بP�!~~~���l�_��Ϻg{��B!�.����v��@����,S1n���3�F�1'W,����A`���˫y�
M ������<�	�Q�p�>��_�) (xx�J���ӳ$@���>�;��G�������u�֋�/�	v=�<��1�Vk�Pr"�ɛI#3Ú
��c��A��{3�TV��]}��b�2�^`�`�^w:�S�!�Ȁ�b[ػw�*��%�����ұk��119�xv��aݳ�o��1����謔���u���td�ͮ3Tݴa� �W^Y�\q�;������j?/�i1i����.�ߘ���C��C��M/��e��FBe�%�]��wwK��;P<׋�vL4�;-�Z螜�LNN���Zuٚ�O�'2�&�2j��RǠ˒��+tԋųl#}�?YE3�*�"g��J���0��\w��d�QE�4�3-�<���㽎���� ���1��үQD,��I^�xD���7ww�����`����+�����y�Ǘ�� F��3G���&R����'�����<�����#}=�'jj	�)(ʱ����=�s�����~�8��/����`�,�����߿^������uN@�@z���������ަ��>L%�GɅ���H�a����=?&���� �Z
��A��M7���5$�"���M3�c�7�K�����Xճ#w׫w�������g�C9A�S9223�+q��)����e�SKvXy���y�R���X���Տu/�t�I��Nv�)7��w�5�ET6OLMi�߭�{���ق�@�^� ��z��n�Clˣ-v�j����D�Au�L���6TՒ!A�w�v�'08�&Pd���ԟ������z"e��W��������WH�+!��<0RS������#��T�Jl>���\�7�y�b\DH��(k2��R������\Y�p�,}��Xчp~1q��`���r*2܈Kz��;�?�[p����-C*�U����F�ѣ� ��,B}���]E����W6�����W8��:����˙V�U~�qz�CW$���8�R��p�A���F[3'��{xyAg()t��N#+�l�n�i�y�:	V�H\�?3�%�_X�tʲ��K��P��D�H��T���GX���zb���?A�|4ԋ��gh������ʆz�����R�V��;1:��E}�����c�L��{qR����@�o(71�7$]g_0>h�I\T-^��2�����NU��˺�˄�>��X��ve؊} vk��ս��v���׃���v�^������H����2��t���Idxz�+˙���V�إL��#�9�+b@0�&m���Y2�����õ������"Ͳ��e���/kɻ�%��|||F����;M g�Zg��Ć����bP� �������Օ 7�g{纎��ɉ�h�W[�ZPPu!=|�Ӗ �<�j7�;1�8fƵëU�+0�@ �A�������&����,B����A��bT@`��Z�����
���<G�5�ji�]�k�Te�XI	si���b���o���;���>_�|���X�P>-!�H��Z:0 @�� t�n�V�4�I_�_��HveH��"< �e.ff��2y�31�˗ek���"#�]�ܸٛ� ~�V��O�Bg'�.n5oX/-L�}����P�2+��44d���_����y���McR-��]�p1h�B�Q@@ /9����� 5zC!���W��iS�s��&ݠ�`2�3�Y�5��Rg�����yp��>x��It�; }`�^�i���< D	��>:JMG6P$y���s��@q�CV�ʖ~�6�,�*��!��|� ��Ə����R�刧�r�����V�M�_#8�!����:N���s���T��N�%O��I�r[����뀧�{���ȖDF�&;������{��%E�B�ɼdeuɸ��[�w������^^�zq���<���>�9��ያ(���9����	bv�����.���Y��ƴ���I�?ƨq����ˊR�,!�}ư���ntH���j��l�ЀO%o�|w��r��ࡊ�
�z P��
��%�r***3�TyU��X�$kR���d6o��pQA���.eP�]VvrϞ�B"�VUz����b�e{t���-̟,ݧd\LJƖL^�;��P�n��	\�;�S�	���_N?� kK�d���nãM�����*|4򶶶�k��J�H��n��DI��j�<i˻��UE�����{�\;'�'���۵KF<�S�8�U4�D4{�}um�_Z�����(oll��M�]RR�u���cecÙ��I��a�PV(ʬ��N	8a-_���`���Ι\1<�8��DO�#?I6�d�cMP�Y�|�Z��_v������ �����"`��
��w�[3�B�w���?���Zy%#��Ձ�m�}S��p	6��^������-�\*��e��W���~*��>��o3���?M���m �-3队��ɛ���c̓�����ۺ������'�\E{|��ŤC�<��`x]�Z�8�:�w�_>*<C��D�1l���dffC�f������!o��@�	�9C�=a���~��v��~��Nxa-����R��"�DU��-��X�Ȏ?�ݚB���CB[�f66���,d- t������������ä��3=0𜈄�P@l���۾� �]�())�'�g�e���+*F���ץ��-���gw�*�H-�|��8�{�oi ���m�h��M��:�3�o�pK�HS�7:��|BB �fU���BV�@�P�p�cT���z+$ �5���^O&ϔ �����|���&��R��n�I}���3T��b���k�2ψ��8FOLL�~k����`@�V��ŎS����p�W�ӳp�@'E@�M�*Zjl[PPPl�y�1-/{ls H��co"b�V�J4��+����Qr�?�7��Ӊ��#E��-}Quub�^^�Y�3g��i��F�Mm��J\zE�0Ktbcb�Ok��t�k�xJ�'�jV\V�����:�4�hċ��N�s���M1�EC��h��|��4ߗ4��:������Y���g�� ���r(��'��Ć����m1�]�`o�����E#��>�tĊ�[����ڀA D
�d�h=�`.H��+.��N���N�&w�ی>���LZ7�L�j�OW[��d]>�,Z���p~@�A�v�|С�Qj��������c�%�ۘ�o"i���㳭N'>|ll,�U�]⌯c�)~�ߍ���H$�R�L���ʀ�? ����c��_���zu�¿T�IV[�rp��@O�gW"[��\ӇƩ��M~I����W��>~�S���a32CZR2��"��Ġ����%+���m�u i�4��8�}�(J,}��C�°N*ᅟ[FǍ�O����*��%GwR��g�!����Px�T��C1[}*  �/*�����\��̗!;	J�)\k�쀑�Y%wG E�!9���2&&�
_ܵ�{H)��^�x���ː4�Z�p63�pF����S��CCG���.o��70`�l�71��u�?P��v|�Zv�r�v��p���f ��d���Ņ߮���fff�f�����-M�<ey������%a��� *���c!8ɺ�������W��&BW�%�OIMx�h���0�S�o����-��-��dM�4����p���t��I3�d�����| _���n�d}�9`G�S�Ȩ}y�%{ �~���/��?E�?A�1�Y<�L�����������Z
|TH��?*�V��*v������ӝVPk��&z�J����1ۮuF�1Cg,��U�N�_5B��a�W�OϮr#���
C��_e� �N�B�KD����Um�M�e��ck��)���悫hE��|�s��*	"^�2'���:%?�wH���H���3�ΐ��/�!�sgVzM�1w���6t���ʹ�P�sW��߿	�^a >ĉNQD��Bľ�Z%�W�G�kU��ځG�05���C�A� ����i�H;�M�l�0����C�]a�/\4����_���������P^� ���j�-9T.
!��J���?��e�.���z����5��
��|h	`�CR7�t>'��K�J�H�w2�Oؒ')�s%}����_��ڎ ��MMM'[|3QP������<Y��e}�rg	 �1�^-|Ipï��jf���F���6�%ե���c�[�[�{�9�`��Ƥ~���Qٜ��N�M��AUU�`��۠$��'���g��fvvx!��ؼ���ۂ:��P}ԗ�@;���$�F��;6�ݵsv��_a�����:���D��zM�C��\QW�T��s�Ez2�7���w��_>}ֶG���a���=Ӑ+��F���&ŹAnD����Z����(�ۻ(Q�ϒ�'*X���+ˋ[ޗt_w(��q��Ͳ�q<@���`(O=��w�僕��S�
�r=AP��G��,�z=�������3w++��^a(e��=(m���J0s܌C��E[�7�&*7<1ƛC����]wO(1���z�Q��X���\E�恢������<������h���F]�@-�N�;<P�g6�P�5��CE�ן���@�+��P�>����I����Ñ���Ҁ N�&�a������nWvΑ�sz���O��{�ePGf��9;99�w:����Cp��0�yĸ����J���G�^ӫ�,d���	hJ[[[U��o���CC.�����:Nx��#�6����OEi�Y�k?z8n�UU�`٤�w���C����Y>�?`W�����~� �c$��3D�v�>���\ʹ�E`�^[. �YZb�.�Rק��,R7��|P�G���qCՈ����1��S��[�7��HZx�<�ZN+m�]
���{�^����H��N��Ъ��j��6��W�ͪLU��Z}j�;������֞��Y�ė{�}�?~�}(���Çe�(Ct�U汹o���R��}뇟���&�)�C����X�Ǧb��w�:[*,*m���7�����Fh͘}��nYqoqn�����[���-O��_x{�iݭdg�m�c%�E��ҳga E�� #>�ֶ
,�K�)�?Gj�i���8��)`P���� *Т��;Vg��,G��M����=��;|am�p���N�L���,^����}�֥P4S!�U��"UP�Vw����d�����/SZ�PrI���=��uI"2K7�/7�mdO����.N�R�.YK����t�[��jc�{�H'�ڴ~{�S9>�I����pW���wxSK�m2^0�R�����/�y@�@����&�y��� ;��jj�������b��H���M��{
\T���ii@O�!�����986���f/�+++��z�Gc�$���\y�Dj���\WwMH�6�r�`MZ��lP���S��	����?B���+<;@LL��9r�G&�B��<��yk�wdd$�����M=��J�5��~�����<76602���Һwс���*R�3H�i^K���O��7���g��}����	�+>11,2���i���j�g!�K\�md�r.���}����?���,0�}es'�#/��k�$n�U�3��QN�e��IQ{�'}|� �9�+�-�c;��v��/�)2�j�2$6�fv9
/�G�C톨�s����t��Γ��L���cy���e2=��F���4<�t� z\T �>��$�}��a�X�|B��c%�K���0�k���������{�j����\\o��#b�?���T ��q�Xۢ��xSX�B�scY.vv�'O"����7"�766D��h.�G��P�a-��O8����m�>.�����iii@��Wp6�캙�sOb��&r�&(i�xA�^t�tX�|ǲ\�O@�uO�
F�s���4�z�M�^�v_	�w����Pў%�4�)�TK�>���$�Y?���Z�>47bZ`�!a��zr_�b���DzNO;���=״��=�����8E�e��P=�[��-,��SoG��1&(������#����/.n���#޷o��&�~~~P9��u��N�EA�hi)O3���<��켼'u��\������;�=@Z�j3��{8���{�gM�ڵlQ���9�<|
�VQk�~����o1���_ėu�� ��E��aqT�}���i�eGh<�E/�E�7�r|�g�ONj��hc�d�N������1��N�rr 6�BKS�ݹ�l���7느��B&-u#���4��w��ئ�Es��o�^�I����B�|[!19y�m�N��s�c~�W9�p�G&n�[��� &����<��M9�v���oO���\�s��`D�Zȴ@+���3���ӵ�P�٪G~/-#:���IC���dA����``@��.h����P�IIX{��w՜EbM�W1�c�VV���;�
�/> �Cԗ��6���KY//!�L#�o(U��q<..hV3�'����o��[��`�)���	"Z2��F<��k�c�¸�F\T�@zL�uTpiq|D��gYæ�����8ێ-K���,��0�RX����
��:����u�������VN��\�p(�)kk˖ᷚBg�r�������獫S�eH{Nr4�6S���;=�����t��OLN� _p.��a˄OO��{�n?UV�����`�Y,)#�����̇_PpY;��?�	�����o����z+�G��ɩ�����M���K���UD�����d�)������[��x�?�J�4<6)��� rz=;(u{��??L]h_B��L�9A�&Q	
	)��[e��W��nS���q/T�e���Y_�਱o�;�Q(FG�����U�r��Cu0
''n�8�	��Q懇�fVV�.��|D�/^<��|���[�8�"Dxxx<����~?	���
�t�j���"]�}`y�.��A�Nlt4�(1@= c_�� ��{���@/��:O�۷��x���X` 6�wuu�"����=��j�SA�(�뗯��b���|Cs���Bn�Y)��=k�Rőy1�>AA
-��p���~
2���
���y����Ƹ,""c�#�f������ͤOS7��	B,�>�m��.!++��~�y��Ox�� {�S�ih�4���ʏ4��N��ΩQ^��*J�k��C^?d�Jr����6���U�{���x���
��m����mz���D)�6�����8���9a\�M�Iٚ�99y�Ӕ0t k_=i��H��t��:�����ibvlGk��}I�{@eCi���P��:���3([��L��SY�Ϻ�Å��7�;{�����tL[�T`Y��O���q'''%v��+��R����7�2��rC�{+��2������������[�K��;#�Je�[��������ݎ*�7)�m���K��m�d8A-���	�� -c6q�5fF�*CC�a���-�$%@�L�:ls�ɰ�f1�ej$V�k���L&�#""�W�q���C��xD�kj,@Ȱ���tfH��v`����Λo��0�hx Zi;f2�����R����i(�2���-zV�Ηɜ3�P���-����5�jޫ�:����ۍ��ǰ,�p�G�Į���Q�w��$�T��hl�FF۞�j�]]���02�����Ƕ(�:��]��#je�� ���/҈���d޻�_J�8]-���)�	~?��g=���b���j�R��lPs��lK/�"�J��^^^P@#`��������ւ�rR�Ҏ��2��Z�A��1/���s�/�1�!y������]�g�bǮF��v-�o7�����&|��(��=��xgG��G�&�W�;v���%ϻ��é�����A'��s~k�������)�d�������n���*Gff�Z���s��W�.�&0+Bլs5�댈STV�<�ͅS���w&O]a����	3�\����`B�
.C�HH�r5q�V��?2��/�q�XT�����l�Z����?�7�J
�Y���.9��K�X^f�a�Jxcjbhxw8uh�=Z�c!�	�uW���x���C�'�_5�K��4�W�RgV&%�-��]f�nO!���X������ӡ����{f?E������Y~�J�Ė�l��z�B9:6��+h�0іێ�~wڷ��H��`����K�(�9h�GӠ3�2��*"���]_�a�w���8����;�|*�s,���[�=�㧍�����pt�G}����/^�9�+u�3.P`\UKZ�x<���りwf�\�m�5K篽�g�vC��]NP��f3:���>Ȅ�uk�������/v���E 6/�O�.1��ȡ�����O�?�_A�'E�P��R�[�\�����^����'$��fd4���l��a��3�Q���IU�R�tz��ۀ�N����c�4��
��9c��,dY��.{��~�)�e�}����3<��ke���_���ᾤxQ*݇;d�غ&~J��%N�=��7�˴8�}�w���u��NӖ�d�wO�Z�%����V��v	i���|-�,s�g	b6Ƹ�{��~'��F��Jv��X\B��Yf%�B�ΥQOY��?*C]���R^W�:	��R��ѧ]v���@�E������`��O������v��X���/��Ѿϯ.��gַ���<����g�Z�ڽ/[����`��߇����kh	�W ������������?�b�$���y���Ї����p�'����k647���.��n�خ��hI�B[��!�}�X4R����Ç��.������8E� �|���T��4.�>�
P8����S�0���׿~���	�r�� �Be7���x{���khh���Ƨ��@�����
�1�t�o;xRSV���	��"Y^�"���P�ָ�"�Z�]c&\\�搱110g!������?��@�҇\�� PC����@��}fVɬ�������A4h�������lu�<Vd�������Th��������ğKH�8�����{�6$�@(<�u�	l���8T���	f�h��ż��aT�U���qpl{���_����c�'"f�9G��s1a6^�f�9��BS�u7UUuuV}�cX΁* �C�T��\���u��im�	
+8ux����^Y�6-�����Թ[wRn�>t��O�Y�L�K���8�麪���x�*����|�Q�k^WW�o_��l]O�(��B�8���#e�^n�Ø��n��-��� �w&�L����i�ZJ�r���h�%}�R��<�.������Ղ�о���X
U4�Ѧ/pg:$5	>��8�<=	��_��1Bw���KK��8��(,*
ډ�&N"}ٿ�c�x�iJ�)�	�z6�fc��e�gPTXxy3�
��tΆ�g�2�8�S�����ܺ;�������A�o~���`���$wG�{GU�c��9��j��KAZ`|���nw���k�J��������ڲ�7���kX׀�y<�	�l}��қ¿5 ؊9�wY�g*1���}�}LG���f�����R�ޯ}S*o(z����S4s�|�,����D�0y־���1�� �q�e%P�?�	���=�I�ǌ��a�t��MW@�}%jܖ���ǚ�qS�%=�g55<Lq����<6�kj���WQQ�-6T[)W�����l�vl�ڀ�����#��-u q��A
&�@�J@���tx�k�Cg���A���~����>11!)�f�ѻ�*AV��[�N�wUX����el�_@`�\Y�<���)�N����3����G�}�AF<�Q�;����+y1���LP��f�b�}5��ȇ�A��7�4�
��'��F���^����N�> X�vqW-]�r��](�lb���i�Y�y����oY�{����>I���`�c@6�F���a���z�S���O�Nfߊ{˿����z4L7Y��E�H��z�Rs9�4�뛛m���B"ͫ3�o�Ն�����gz�z�[xa�z� ���E��&(o�6T~������tk(c�$	�G��\�����������FF<Ӏw
@p�c&9�j�8�y�@���Iu%���7<��葲��5z7S�~����A�uL��-��޼l�Y��qm��j�����lÚG\"�� Hggg�q��>zeb�����n��| kT�+�,f ���"%��+�R��3\��?]���b1YY�@����פ��!���J������v}�����a���]��s����*]	������q�u7����G ��+��l�f�r9�L���Oɏ|+**��TB-�|�ԍ;��~��G@�i�:��Н^��MP�SۘC96&�6�;�i�͆.�B�Kj�Rq����=��1�XqC��Z��h���w2�1���?�$yC�Ws��A�f?C�f��s?���U��a�d7�w괹y��`7k����!\��L8��l������g��)*�@�/���W��r�)�A�I�ξǩ		�4D71�uJ����j���zM�us]8��n�	�Rޓ+<~/&��d�$`[�WR�V�rs�վ�2���i��bgi�J:�Ѽ�}�uľq'Q�EIE�ȏ���"���OA�kqoT�$�dt�&\�wo��'=<�x���w�d��-\RE������E(����
������^tDJ�$�C�oP֪�񮈥��(��v Vяʴ�\�L�w�8޼ ���:K�(k��L�6�X�O�����"`�0�My�|@�iii/w&�о�����t�������P��Iq1m����o�C;�����?o��nØ�ynB9�@� �u�q��П�a�-��瓻BM���q�-���#��R��*�ʏ%�ܻ��̹��|�B�O�=�Ul�=�H���sH��#���qiii�N�$ǌg	�� Ul_�<#�i% ���)4�N,.Z�1�h-3���
����Y��	����N���/!�j�L���)|�}t(f�1A�I�D����PYw��Ǿ����� �ޢz����S���u�"t�r���q�X�F����3}==���)�	���X���ѩ�����"E�j�D0�Q�js���<+��V�u�~�2#���x��"���[�聿_�U�obH�|c��sc�_@����
��(��Y��%2���[�u;
��� ���4�����E��G8�<��	�p�^���S{�4�4�碂W�4��z��>�Ot#Z^`��}*82.���ɶ����K[��ۀ�d��Ц�Dݞ�&���Y�ʦ�����)i�wyI���sch��Qn���_�뇕m;�nW��^\R��[D���7/�4���	i�x����/,,�� m����rA=���-�R���o^#���J�Xx!S->jd�����))]8S��)]q��-*㉂B�.� ��B`o*�]�k���(o�{��}���Hg'�Z��>5uu$�嫞��z\TԬ�1�A��<P˯���C�C�6�-X�V�M%�r��������<���IP2T��9X��E(���y@W]]}�U��iL*�������V�U�*�% j''�k4<[�Y�	}�+d�K��c�?ZϠ_��|u�G��7μ]1�lgq��;zI�;kY��n�qc�8��(�"-=��댠S�9V2��>"F"�w��鮆��~��)���s�ۯ��===]��F'.|����M ��A�,���!��9�---������������A:<�k����[��9��rN=��H2����o���6�L	k-��ݠom�m��]XR�:?�F��m%��%-�%w`j�a�uֈ�xc�V!�?�˪�-3�uMM�ö�m�����%�t�Aɻ=<�5N��&�ۺEkΈ��u2v�d%�������r���U��]U����ؾ����&1E�?����?(?�� ��9�������B�^4�[�kb�|�6��e�}{@5\O�·���'],���ۼ�w��5�8�f���jW���XP�� �PLdr�u��B�*1!��!dz3�~��Ն�T�cy�%�]�ӛ��[[����]��fi�H��W�-$�C�~VΥ?U2��E��(��P-��Y	ܑg"����r������0n�$��B�%W�����T&	b
PR�ʉ����@"�ZgwX��XƂ..�����ikks�vw'�u�V%�ʿ=�޴
�/�cF}�M���X���)�A*�~H��,�{���YZo�	U��ׁ��ԧ����?s�������rl��c![�[�8г�eg�	������צ����	�:W�"ɀ|�۰�&��w�i�7�0H����@�]�7u�l~@YY444{,ۜ�6�w�]5�)<<L���05L�& ���l�������u��9�&y��(@6��bD{T )�HV��n'@���0ܹm�OeG�n{Cɛ������rs���-�ڷ+J�:�V�tmx*|ew�4'����N�ɽcrX6�L��/����� m�w8��;�hr�b�M�?#��%�"��V�r��> !_����tkILX8
�Re�.sR�F��$w����R[���Y�変��z���^3��L/H��a�6��Y�#�E��U� �3��3jo9G�ɡ8K0?Q����x���{o��0��zIQQ�JWOO
`x�%����Kٱ<�S�A��Q7����YBe��X[[�\[?:�=�G�*��]'�ƾ+��g�g��!p�
��55눡4�\xEX��k�g��C]E�_wK���9˝����e3�{&�5fii�y!��}����Y�/AMI��sԌ3|Ϯ3����R���[��Mh�h~!�A��ܼ8�l�Ǐ{��O.Źm�_�ξ���xM=ō�&�U�n��גּs�H(����O�>������
X�a�'��"jsM	�����G������F�>@p77tCQ/����J��Sc�ϰX�����X���456�t�m?���������2�9�j%%QM��98�N//�x�LGC�H$�d�6�C*ݹ�h4_����wh���~�L��*�Hz�W[��6z��xkb�cN:���d7S�F�w��6�ff������TSW��^>tO�������h/+��c+���Y�]��4�
�Odc;, װ��2;�3���!Џ�n�>�=(���Ⱦ &�j	]�w�����"�N޶d� J�ym�����Ĥ�}*�su|��R!7���x}�%#�}xJ@JSӮ~Fշ�Bz�m#�v�W��%��� r�c��#�O|�A�!f���>/�����|q�	�yxddʃ�:��2@�L
�<�H�އv�����٥Ζ�Zߍ"�G���Q����؝�Hs�`��iޛ�����A�<��+����7��st[�|W�W.>��� �5^�_�!��j�����1-���ۥ�TY��uG�V�������uXj�f��A�VV�m��������͛7G�8|VG�K������Q�A㡾(헐��so�7�i_�#�z����Ɠ'O��գ�����*���e#K@�L����6]@r ;^��]�A�r�{��Ԗ��5�Y�'`��P���k}�K��>��K�.�J�4��צN��blgoo�Fm(a����(B�x&�����1~]Դ8s���D�A_�3UU�p8�?n,��jR}�����w3���/D{k��K����@��]܈2dd�p"[�R��*(�~���j����Pή3>8�ژ��k�B��9�k�u��5�ޭ�*���\dֱ<������	���_tO-#���s�Օ=_^�*���|<�l~�qxX2\b:�v�,���-�Q��Q@�� �	�N�Oy�g�9�B{��,��f2At	0�uK���'$&�����=}�t��N%�o{��R�4vyMM�����	J�k+++Y997�bp,����4*��x��0�� 'ww`9�5n/Jv�e���H���R�ک�  ��rB"oޝ��,��7y67%i��V6N�G�]LȿD������`q.D/.��}G�~&B�ԥ#
��R���+�G�-3��\��H�"������m3i�ig����_��|;�!�c�v��E'����h_��_�ť�*�|�R�X�Ku����^ɬ����('55b�G��n:˦�c�xU
�1����`��o߾�$��cA=��m�����ض����P9��?Oнm��ʙUNB.e}��Y�
��=ܰ���s��jppp��]�ϼ����4�[�-�x�q;��v흗����a)��Sv��o�x@8�o|m�>BI,ypU�kgrq��)�Ǌ�@�>��si�&�eݾs�N���05�w�������Q4BCO�΀c�g��������*S�ܜQ��ۨ��;�Ʒ
�ɯ������I	��R|�|�xdX�� ��O�=#����3=V"#�8m�n���-���adlYZ�H�6���q�&V�9�6����}(c
c�a�P\Rr��g���`�PgF\�-BކС<uE_�̩:�Ҧ�?����<������I�S��  �Z\��Od>>��Qp�wUݱ(D� ��ۋ���7׉��	Q�p+�$��+�*��o+�ݺM�lll$�=��� NPj�!����OJm��S��Ւ��n��M�����eKfL���=	x�����)Cdddk�	L�*_��T�PP)w�ˍC���t���|�,x�}�
�?��"-O�gb�[��ֻ�����R���Չ��F
��V&C��r�+-cX`�l7�>uj�S@�Y�VoUFQ1J�pڄ��ŝ1����
��pZ�y��ׯ��;��4*��&n�8�C�G���j�4��],�������I6�ލ�mz#2w�1�z��H8S2w��up�ƭ�v:��@_R�^�e@*����&��>44�6a��b'�O�!J�_: �J$��/D��wW�ފ��( (O�>;{�	��%��ĮڿP��ϟi�Y�������`X�Ӥ����Au:�OHU�b��L�


�w;7<��z��?�Lr��	��ܫ8�&��f�nt32�44��:솉N�8�	���*��G)��n#�近�t&0�z����6c',���\L�=)������ �j=� �����TUQ �3(���%��_noo��q ��^'�|� ���x�,R!g�\p�b�j�|nv�<N�RlWs7��@2������@=�/���p�f����Kdfu���J������ʪA�m[��˄禰������f�~���\.�)����!H�g�r��>.V��+)��|��g�S�Ϻ�l=���f~P>�	~P��U�J�e���t�-�ݟ�/�{P^��:���������R��W��-�h��2�����O��>u��<'S7P�4� �9��8��TTT�\��I�',dY���rDo�����46�p>{ <�z�m�%W���i��s!��c�n��%�WDm�}O��Z��svjiۘ�\{�>�5qᐳ�J=��5'-N��hW�%X#Tm���o��RQ����:	�q��immEb׏�oWT�G���6�n/�� y�����`,�^��$n�H�0�K�muu�����-���Xs��<�WaŶ�6��}C�A-U$�<��-�D�Af2�N�tPv�����˅{����K��$%�5�3���+��L�IO<q���!0�v��*	گ��x��~�1��f�������?�ڍN5�?�����pm0���8MI`�g׿�[4򇴡=F��,X���ʄ�4���@ ��q��<�����
%C_F�
� ����k_[o�+��n�Du��mj�C-���+D��~�1�F����/��A���ڋ�S��װ�g�t�H7'+�q׽� ���GuF�������QdL뽝�G4ccb���H"�*܊��H�;na�ޅ�,:�z����Ɵ�n/�Ls���BK��|�8H�O�㥟�)W7tZ��LX�	`��޾��ڴG���o� jj���.�1`�����x��������k��b-*f��RiоP+�i0Z�k�:#����\� |��[�ÖX>�ţIς^�3��&ֶUp_m���^B2K�
����1@ȵ�)##����i.#��o�1m�k��r���~y��j(��tlΕy��$ �!�%*�t3�Ž��OY������k?���w������n^������K]��7�0t;;< 9��U�())A\&9�`ʟ��߾ڨ\rv��17�����R�����>�p���oPV�IX�S� ǀ���K��)�%������+Mww��E��6i��F��iO:P����:e&�3ɩ����� �a�����j.\� �`Ȣ��8_^T3kxl��
�8�Z����\������\E�u�2n����߉�?��"p,���Ë��s�&�DXX�?��e�"�ЬʠD���n����n�J�ʪ��ꃮ/����R�n&JA'(�����n<}�q�b��ؑ�Մ����gޡ��7��R{׷�;~���4@�S�X<d��m�/v�W�����ᓓ�A�#�B@�7�
����wS��W�˶.��W��.π�Jȋ�U<`���.����<U�K�_�7D,K�xƅ{���,)�ZF���߽#�#�0��	�=\������L����?*c@�����ʧ�EO��,�]*S`����������AI@3�+������Q*�Mn*B�{�ዋV��rL	?��۬��^]]��Su5l�"<��Lxt4~�ȟڲZu�,
�TS8�B���������{	�>����sI��D���ȕ��ݿ� �>����'���L�o	@���4���;���T�"�<���;�\��a��+֯�����75O�������zM�cT~�칞�h�#~T�+0+���3�>���/�%���%���`���ɉ��gx����h��'�>�(�3���@z�f�O��8�b�kk��%w�He��;wZ8:�:Rz�����8j'(�{�q<��낭X�H@��	�������F�aZ슆�&����ToQk9߿�|�ä���]9K˜9��i��Ix|������¯����=���I<	�jTMM�w�D�_�ͧ�;�����x)������J�L:

	A{���������ڟ�ݼa`h�id�q�Hӧ�:�@K��������_Q�Ga�\2�������Zyǫ��GE���}�"�%}{B���0@�����W/��H�2���l,�oy�5!��v��{�NAEuSbu�%�v%ɰ5�)A)�`��JʹR��7�_7^���
�߳��e���G=�9�(��YNT�0̠{w�^�������A[���H ���

g74L[R~��'"&v�t��{yrG�U��o��2�E�I�m�/��&*���f���q.m�k�� ��''aM|�M*����h0��ѣ����%ؐ���i%Ќ�%�It��r��G���������Z&�w�{Ϸ�H�]̇U�k��9���Wf[��t���k$W�9� -��G��aJFw������4䕕	N�t��x4hsP�p?���*v���OX�j���Arw�7U��"?fz�e����PA~��"�֑\Ј^�K���<kKAM큸u�x�U�� �f�Om��b�>�c,/�"��)~�Fc-���( (�qF���ݎ�WRQ���a% $�j�Ɛ��<�\]X�"���ۿW{!WR�أ7�L�8��gA�Y1V���%M?fv>�Hf�i�ُp g�.�␬���$pn`gg�ҖQD1f)*�@'�/\|>�����_�x�h�˕1��ѣG;1s�0)�����!�p:F2�mJb��EA�g�$�`����a��>ЉQmp��@�ល���cKKKR�[)eYYY��J�HHw��06���a@�՚�� ^���e���Ϙ �Ҭڠ��P_h?E<��TWW�\'�}Z���NVV,˻�\ݭv��t()���C
-m��hr�0����O���.�;�Z���jJ��pW�t7��1���؍�/��]���N;x���[#o݅�#�N�Y@�.,*��$"c3	R)c�C�e"o�<zerC��}�<S�k�O2���z���s;Ĕ\!�Í7��`Y�ww�gw�S;,^)���J�w�,��E�$���='(���%�Z���kw�-$?���3���bs|�h4���\T���N��"�7�H9�ɴ"ϾC4�js}��9��@�m�ҳE�r���+���:��=}@˵}SfI�y^�,���k��p�]i[�Ĥ/X�*������J�ѵܯ_}�����ɿx�B������NÐ*�q\� �`�F�;!�u `yCuV����d�<�o\&��|ֺ�۱O���"�-�n64H �i�k%�Mu��?�p�<�i�]=��eN
 �O2�6��M��.u���\o�6��W 7)~b�4'�� 1L�T�D�q½|	g����k[�;�5P��woOԄJCTUa� 95l/�pOOO�WML�x�jj���'�@Y	

�N���Lx��+��|�~ivu~d�r�ӣ�8]Kztt$����ʂ�<S�|�⡾�a�d�q��k���Ol��n� ��鰀�m�Jy�3��NQ{���:wySHH�<��S�:�׎�'��~����G@i�@p�ڠ��2��+p����`��' @���s�t��x���∐�?��
|�Dg�!!!!?.��kiiI�{���������###vvv{J�x��XI�I���Cy�]L�3��:�!�����{��w�^R���t�sHu�1@��n��c���6�o,�� �"�ʝ.ƺ-��7?a`ce� �y�;������L�I��E�7#���o�"�O{:;쟛#��.h ̅S��M>�Ԥ��]���]���O�:�(������ 
yU݊&y�r��H��ڌJ� ���c�7�^��\����n̿�n�y��s��]ZT�;Q��� ���ǘ��M���������B�N��2<f47���d�]>�]�b�|���3���"�MTK�X�ȫI�ɀb:��=��0o����P�i*�b8LJ��v���5+׃�Q�a�󫽩##�yHcmw2��� �e�U9ͽ{9��_�x��Ƅ��w��Srlw
S+("N.��O�d���5�7��gƋ�R��O����f�L�B����"�_?g1^�G��/O����z�}_�u�����FKK+��
��UUE���ӿ�	�e|���Բ]���/$�y��}1��5~�/ss;v�oÔ?� �V�5��	��(��F0�Ƴ�-���N�J9���1~�M �j׳ck�ʃ� �_9�|�k�0|�ޮ_È}�Z^����C�*kш=`8G����ݒ��"�����]V��@��,&".�Z�����PU=_����DD��P��.��R�S�[�������������Z�z/�̙���93{���\�(Q���Rz�c���0a77�����x�㎺48Ȁ$��T���IS�����o>Ck5O�vm��)-��(����g��.)eff��#���c���������2_����<��968� L�(�^�y���a*�k/��U���p��p��qqp^`!�������k\���;�z��84�ZT�C񇫐����f����%@	�\[ߴ��M�zz�f������+�����0<��d��Э���|�"*}�m���aRE1d�w�����nxr�k_�>��d�W���A䅯����傞������zK�|�dA�(�dA��oco{��!JZ� d��A&���%���e_�g ��jj�jj�NvP�����T��j��������/Z�:��ڔ�����'�ŅtXeMP`M�������AiU
�T
�Lv����oӲF��j�Ѭę���85���D��22`BWm����$��R�c�^KA[h�ϡ|��U~�]^����P���JR�t���8f�غj�)���X�ҩnW��3|�M��y����7��HfSQ�����o�z6l�44֠���6=��c;�I-P�U'�j2������|#�:wu��j_����f���@�W�x��΅����41;�A�s5� S�x��H�"+'��?r�R��z���u���<�?����=�A�|��gG@�e�&����N�Ƈh���?{��k?'�����v|U
Cϕ�+�"�����58�c�X��Fp�|A��:�a2D��ԏ��G��B��#�WNOO�%�����|�|KB�/���ȣa\�����[Zh�Y5�I�5���a��2c�E��e���rV����3�ű��|��bvb�h��&�����Z����	�'���ֿ�"�IwW�Ъ� @���	>|�| ��Y���\�a��c�'gҹ*.���֖bT�,ϩ��0��̀8X�S�o�����j�:=��?�iJc��#��X/�-��,�װ��[{s=�̈́z�
���������M�$�%�S�1Q�7���Ǐ��K
�>r��2���"�32e�������֌+p�������7�2	�y]����KuJ�J>T"@�(�>䨘��F$�����
O�W_u=�-���q^�A����"gg��ow��l�&RI�+TX�7��K�A������}& ����"�ST������%��b9S���������G�{~^Z�9>p�B�Q��	 ����D��9??�S�a��"�{�4����̈́�,�b��}GH8`�t�
����)7讛KLL<��W2JW����"%��$�vz���GW6U�m�������(��~�e:	99ƿ��-h?1y� %�&�� �R����'��2�Scȍ�팁�b!e	�4
B642ZYz�_����i
��%�~�7SyuQ��7���`�~���%�=�F������}�&���*`�9�|����|#� ��M�&��>)F��r��m;$p)̀���2��;8���p����R6&T��ZĦ�y�q�%�(�Ȉ��D��\�"E!�� �(iyy	��������Rε�V�d�72�����Ы�)&���Ã&f ���o�>��y;L��"]}KK4�z~�ۑ0I�_�̎��~ �$7�F�T��X5����ԃ��t�ྫ������+Zy��ď@�����U��5E���̐�[kJ�}��rn��	����R�h��%��{�U/]�.j���\�16].��w�S��;���X7�1U��.9-yp��� S�L�ͅ�6��-()�TP� l�Y��uȯ_,P���~C��7S��''�%-�
��^�n�[��T"
VPT�}i,����Y��sT������T ?�DyErB�-�ZȘ�P�.:�/_�u/E��� ������S�\���(%��s�o�ao��Bg�h��@�'��������9�/�6>���]I���<���s�إ���0y5�u�L�[��O�1r����lܫ����*s \�
#�n6��e�y�Ԫ�
� �,M����9>�˳mh�S�+[Q�2�E,+Z�&�SӞ���<��rss)S3��]��o��.m�\ _�W!-#�x*�+Ha��I�H��}`��	8�<K��	[�y�qe's6�Kt0Ґw�L�����LOlf&%�q��d�m�EHD��x��%%�?FIM�����������]��k:���>��"Q>�߀�by}�`h����UuT�M��DB�6��S2��V�np�\TTT�?����>�#k���y�����k}��X�w��!+_����i{S�/�����U�(`��Q� �h��(���b3��̀s�~�l骋�85��hp{�����?U�ix�\�����B�%1 �М�	1�9qȶ� V��k�� ��mlء]Q�����E퍀K{��/M��q������}A��﩮��C����A�Z%T����Z0"]ӰAC��aqn��ֺ�Ճ���#�2��S�r����i�;2�xM��H�v���[�TD ��������;-�
�T��L늃<`H;�.el��4l>u.P��!$�ҶC_t�"�����@�(���y�©q�!��W����=�N%C�������@�wcB0�ɉ�"�����MR[� ~�� ��O���;8��|��I��"����QK+sl��3�w�چh1U���$�7�!�gw�^ɵ:[�d"��{����p�F��x����0i�!�a�s��������n"��.�.]��.G%���q�����]�o'��ˇ�]���G�B۠�$=;&=����yX
\�!�U?̓���������Ѣ�oz����J,#�!Ĩ?4d������[5��d~��g����}�m��W�����7���C̊����NW�S�{����Ǝ֎����6UC"�kh�g~"�#��	�E.��͈�b�jу�1�MA׏���M�h��%�$]##���!�q�Q���;^�h�Y��Y��3�$M�#�A�"�)��j;�����^�_�vQ�|�~�p}-Qpy��}���K��]��T؝���ٴ�rneF^"�A��|ù����?��eWc�;��u�2����y��YYY��qy�=�0��[_7\__�Ui[\$?888:=���<�ݦ�
X�l�_��M�]��7[��7���0S�q��Q�x�{vF/����"2���k-##��G�
���q�a��P�X������xy�jL�������`�Y��;���aM�����w}"�A������r�{��+t
)�U���ھ�#t�,̙&��^���T/�HdU�Q:*���@��@���'��4Ʋ��Ӻ�#��f��/��n.��/�C&�+���¾}��������Q�-d�l�>�7��'�����	T���Ʒ�F��B�HB�p[���p�Ğ��Y��|x0V��%���G�V�Pj-aL��'��K� (�� �Z[Y]�lN�|v4YV�f(G��GQ4��1AR���V��\�h����6~If�wd��o�ޔt;�,FL�����.Վ���=��]��|��3�#�3c��z�%_��H������~����W�	8�~������f,X]���˒�G��WUS=Of[�	``U�klH������M��>ⶼ;�I�5�p,�M��|�-�}�@�^ʓ_;���n(RR�g#��a�O106��g��=�yd d]i2�cዶv��["0��R��B�O+*��7-�����^���#Q&�pUK��!s�l�a��	�Gy��M�×�����Y�?4���m�N{���I��@c>0p��ѓ�DErw�ȈNM��A��_.�o�~HIҮ��:��iVY�ת���g/ B�M7h~0	�q�M=�� ���	j��S6/�1v50�v�Na�ЦٿH'��e�8L���*�F�;v�Fhzw{9V]&����O��׽i�E��Gq�'��]+���K1���^":���婼�X�/��th�����J���aO2X�M[y7M�w�A����Hnw{i$��T��.v�[A��4�z��F�ƾ���x00��qu������GO��AV1��G)墉:���������pED6�Խ���ͅ�#��� �h�n~���"��ӡ���P�R�J����9��C03-�3,Sᄬ�Ń��@���%�)if��a�Mx��i���g��$Kf��9��PPYM19l��^�'r�7����E��g�_�!D�;k�U�R%��6z4��6��po�]�=L�aK��f��s��lwO$��Mƀ_�"��+�w��=v�5�n$��m&� �����F�����Q�������XP��]V��q֊��l��%��l�Bv �ڼ�Q�����U^������9zHQ�ϊԘ��
�ZZZ��˳I{gY��^v����3(�h�@�s��Ku/20����#�9�<uVh��a˭�[7o�sm���$`�bz�2MSǙ8>o��M91ߥ���uo�$h1���,��_���& H���ȥ���^YS&��rx{Vn`qc0$?��&�@�GY��w�c�u�r��^A��U��
[��F��t�e���^=c��R=����'�����x1��Kpq�Ia�[�iԾ�\F��sN;�l�G�d���V�u|�ɵ�4�tJ'�[Ģ�WT���m5���8�u�4C9^��E�Q����gj\v�*H�]�*-�� ��wFJd�㯔�>�f���9�u�I��3:�g���Ζ������ci~k%������b�T_�8�������K&��#I��&�,��{{�뛛?f�)��o9r��B>��<U��EE��xZ����dh����^�ٿ�Dw�xd�qrrr�&5M��MTĵ8���裀��D�9rwG5߄�]��3�_ul>N6W���_���Pݐ�v�=S��R�'�G�3e�Fi�������*�!Q��ki�h^�������~�Z[���c��(�K�p�C6���sb�%�E٬,ܨti���ʷ5���F�r�+����.&v1�7�mޡ|K�����"q�oo�U7lZtX��� �%En����1�t}C��k~~>53��6gw�G��y�ݪcʢ3v��O�zQ���&���x�x�
�.����B��;�����c��V�ӯTx��W��6.R��Jά��Ɣ]�ؾHu��'���W	�s�'cg,$R�NZ�3,�h0��s�-����w��/�+�J�q��p�'�y���z��%�0Z`���Z�,3ā昴7�������Oe�Tt7o��G��V�q�J���2���7���ee���ճ.7�_����� gs�E����7�?��#B���q��-��	vJ�z�ԭ�F��҃�������=B�2Fon�?5ge���HL4xU�F"�a�{�LO�؂���3�<#��C�W%,�K��G��.o�����f��+�fJ��2Sk���πw���x��'�t?���ON�)l�xR-�����~�nל��C���~�Oc���k������N�SsM��pI֋6�M��Vw+�X�G�|j�wvȒ�y���T��K���z��K�?90����_����lI����ʥ:&ߏQF��T�[�7ܡ�D�>�g�^�&&&4t��O1��}G�������>�te�X�臐�����|"�d�����%�w�İ�@o�L7q�/�S%����ْaY<�O�}������~���"��7�z����TD�	���j��H�hS,����ˮS���3��8��Vb�o�H����X��5�P�O��<��z���m���h���r�����}���t�q�$]�K�&mU�������8��fgF�B.��k\W�-�=>����al[���g��L�Ǉ�~������d^tБ�[����}3��Z�+��M׼�>����-����Gi��[�S�m�x�^H��>�4��|�{��S�\ht3:))8��������a� �[���Q%m�P��V.���H�ׅ���OR��bݒ��1t�Fo�<&z�;ߝ2:��<n+�����u.���Na��M����}�!�n���ۻZ\\,�,�
��K��ϯ�)
�B�W�&�����`�77w�ϴ�=��6GggoH��lk�o�*͘w�5Q���j�ˆ�����co}g��ϣ��c�Y���mB�ˠLb�p#��j���ձ�\����������Zggg�_�q�LW�={��o�}S��������5�����T��ɓ'��Ъ��9E7���(���FEGkt:��t�U�:�/JJJB�/����ޮ��̈�KHH��1k|]���^����'9W�O�/6�1j'����T�*�Q�U;��IƋ���?�g��B��㣖��B����h����X~`h�%�ǰ��7���[�w�2������!r:���$<Xj-��QZ����K����=���Bc�H��n��Z�P�|�[��F�5�_���zܰ��Lƥ�޿k�����**8����w�k��ag�s�|N�_����^��������~j�M��AF� }Ť�5Z��Ns���Н�ҋ�����y���XF[999A�oq<A�w��y:�wwo�����^;h*���6++��d�|��#�wȆ��r��|�i��t@����c� �7���w�ߊ4J��qC�n�梊��*�+�����v�`}KH �z~���e��kE��y�����C���%EΒ�����)���^$M~k5���sO$���췐T׋� ������m6��3bA�?��&z8y�_~���FRh���	����!�iq��6�r���P%���h;7���f�;���;���~q}}J`_�HHBzz�S=>�<�ӽx���ٝ,������������n�C�7�w���㵑&���k�;������P���r���Iϩ��B����ӭ�嶧�S��Ħ+��-@��%kW8Y�g���W�,g;c� ��m����DS���J����涶�3^���jT�̨N����Ϡ��{��HI�&��3A!!#���*���O��d�����@�@�K����!%~kYP�V��7������ݦ��?��(�[W'gg;�P�Qh�K��"6�Oj��'rh��X...Tn��'��Ç�SG�w(k;;A�v[���3��О�Ga���o��7αY	�(����W���ݠ�_�������+��t���-��!�uG��{���՟&@�!l�gb �p4���We�:P���\}��pw�nhl���_g��Q�]����k��Lڳ��O�m$�M>�?͞9~��Z���R�F���K��	5m�[nY��
���71A�����'�^� �ǰ_n��y��l���]�!N4~�?~�_��R���]��v'ԋ����a���б1��$ev[
�WІ�@�1�ab`Ў� 

�������T=Mo/���Γ�Z.��Y4�C�wFs՚�j�(o!�fp�����s�~XT�'|s�o�v#NJyqqA�����'W���7r �K�Ϗ���
��-��#�-��)�0^
ll}5r��{�m	�r��>�y� �L�xޘ��Z�`�T��T2���a�DH(�5��z��<���Fs�rR��	�Lֺ�|׸g���܈�X)}�%$�=n���8�H��x�W*tw�}� �D�-�uf5��|5&=��T�ǻ��Z�n���%i��5d|�j���� %r�<n���xxy��V�o�ٵ ԕ�y"�F#�1?����C�B��;"���x���̇����̗Z<$g�XXh�#��/��Y�n�c��|�H��B�n���u��9fcy��6��R�Ku�^78*�~��,�U��2?E��"%Sÿ���z���a�l����;a�#R;��&�H<�"(�� �e�ڑһJ�ɲa&6a @�JdH��d`�������3��ۛ������<����S�}̓O�y ����<<��xLr�����jھ�@l����0.��T��!�:"�5 L�|���]x��W^^����U%�pe�]J��Ze:"zB������02>G�}eO9i�W��J���z��tk��g�1�t2�66��"ȣ xI���W'�|�4�<��W5!n����GO�kfx||���J��ut��29�r)��xew�&�A��/���ƏY�����NW[�3<�"ۧ�g�!��I7��!	��Ƭ�	�>�(��QdV�ٔ 4"���!#"������M���o,?����i-�a���!��~�[D��=]��!����t��@S��ii���1[��� (���PL|G��&���Gy'^=��d��=�{�Oͮq@T�Z����~�!#���0:6&aF.�:��؋�3X	4��Vհ��p�î��{[ �o[	H�ss��^gj)�*U���Qv�S�G�H�e4x�O���7�2@?��	�V�V}�;@�k�@��= �d��2��7f���R��7����;���DFb�|
���OቩXY_BD�OFZ�E<�'�jj�w	A�������x���d����h<ł����O�|�n��$Ϫܞ�%jܟ@� FFI�P��1��沲Hqq�H��ع*����6~���`��E�^^�i����a|�}qP��!�X���ó~�ѷ"���M�� dT�U����*|��B�ו'222؝���������P���F`
O��Qakph�d���.�ᖟyK�4?��;��~v��^WW����']QYY(k�k�)�N�R{ *�ONpf����=�*�2��!�%���tT�P@�M�^�q_I���zG�Q4a8��Zi]s���lc"�+��3�&�G�1�*|�1SaD��Ml(1g0�N�f666�9�I�RF��W���t�T4��f$��QL�tt�K�"���~�E@#���{!w��FQ@z�}���Є�K/mj�@�֒0Q��-��^������x�& ���ʆ�e���hh4666Yo�]u|�PR��<��\K��������uɾo3T$MܳЩHW�btLL�i �L��ϓ^�$^��ùZ6���N? ���D�H�����)r�
��Ĺh]5��bGG��������6 �輝x�oX/���I��O��ދ��¦�	�խ-��G�mFF�$`�^�4�p@5��zc�C,�P� tD�ꕿ�}7���c,O��'��gѮ���������9��F�vy@{�9@�%=#��۸ۺ�������Iv�4e]B�V�W�>��<��@Nj��prqi؎[-48��	�?E@{��z��j#n�dql�̻w9�c�) ��5�����K���_1@2 �>���"#!ed�[���g�<��u<T�A�h��H=<x��L����c��U8��z/��ʊ,H խ�4�����+ռw����Jv�߿g�JNJ�i�<37'7�Wk�������Ll�Y ����w�U@��6:�'dK\�𻨌�@5�
*b��h�D@�_.�gff^�MoF4+<�r�u�L�4��Dv�B`7�Z[[~�Ɗw��`��@ᙁ�����"#k%#S�$22::�X -�*DLr<�����c��*|����C��̡s��|�=wWL|����|����t��S	t�W��3����0)���w9�5C�9��ob"L���3a�u�KIKŌ�'uhzD�Sp��*ъ�^%&��0��iu��L��ٍL��A
A��҅�~k0d����g=ی݀�rV@�g�d�u6�u�� &y՟��P��^H_��U�)�1f����RN Ê�'*���v�k�V���=S��듍�X�La]Ȼ���F����i'�LAQmt�RY�U�'�d��cq���W�U[R�J�ÓX��(7�]�%�n��bg�j������5�-�[@,P�Iqw�Jc1
Y��G�!��ss1@-����kJ~cݶ{�� L���� s�iWʔ�OE�Ĥ��'�N=S^�C�	�Jԇ���E5[]Y
b���E5n+֔h�n:<��|E��W�ߤ����y�=-8�y�P��r��Tx
.k�dEԧŨ�y�8��ȵT����X5�_e1��v���K�)18���}}!�<��(�*����|���I��dde�������Us�{�Pseok���?�~�G��VO���̧�1*+*�Sy�mJu[:'�}���
>d�+�p�,���m��'1���������'�AbPM[�~���N$��������2�|�J�4��v@ܼ�����b�ۖK-�Yd�cc1W��r]�Qa�{31(�x�s��3fs5�b�����U��"W:TmTUT�J��,�
՘F,ٙ��`�iD=n��?���(��K�y�H��SV5U���0-8��UԾ���呔I�|�N�N�)sP��a-�_1i^�jjhh�<Ҭ,U/�@��\h������&��8�S�Q��r.�҅"��t+��J�<���X�@����d=�;	(���#�H�W +$PC��8� K��XT`��k
#~��O�@���p���y�tީ�N��<�t�ݙJz��̙��0��o:���i99�?������)�S�fBz:�z��f7'��6D��SD���%O�J����[@
�+�L��-����~@>Y�wvv�O���U~���C��P��x�Z�d��E�Fix` R�ŬE��@J،��9�$ H�8ދ3��M���/Ml�i�+gK&pY��<�X ���Gcw���z��RKH�p(&�K�L�����>gkjj*6)�E9��E�
�,,��ZwF�>nW���o���=O����k�}��611��מ��� �$��\������}r��?�\���v���Q��ŵ�?�&����a��&�!�i��?K-3��@����p8���g��>�8-y m��9m��Ag���R�)���u������;��#�*�	YiiaO�C�>z� �������6�_a<F���8D*4 #����짹U����@�-J��y[Ɔ�>"������B���#��]����6|ōG[Y�W�>��%ҙ3L艩<��H�]A�h���SS�e;�F�P���:zg���+�w�FG�1BJ_��hڬ	6���μҷ�(��A��p{; ��2%/|`D&�'��� `�h`P��%��Og�3�n�����O<ov�4t=h��Vd���f�#��,HG����xnL�������Z�P�h�\����,�>ޗJh�X���Ӹ�6��=EP�mPG�����aR`�~�Q�,1wxG_<�h3�ׯ_���r�뉢��� Zg�m�45�q����x�[���(�|�2:�����w��q?�)����#�JT��d�=�����;bl "OPHH��B���D-���D>>�0ɒ N� x�W֋�3*X'����5J����� �,��W!�5�T8i�lr�p^�0�cv�C�8��љz��ɒN��٭�~��/��[A���g�1I�nwm�ڬu趶?S�r���F����-�̓�?=mm_o\��q��]�:^��A��t�WQ'j3��[M$����w���|��:�񳜁HΝw�������P�G+��/��|�KE�����^{���cV�M<O�<ys�|`h�ޖ���8<�.�f���n�����p� ��4Qt�p~���SH5-1����	�F�������� G).��#�����F�|T��<OxH��k��7���/)�+Z�Z�Ko!��qiʃ;@KC5Š�c Z���>~$v�<��
�jv���c�V~��[{w�T%TU\��ZWX�ݖ��Ŝ���)P	<�ׁ	���h���U{�j>�:c=��ҡ 4ΜYe`(�kG�ʾ_�V+�8a�f^��o�BF����4��D'��,�B�lx �9��{������,&E	xu��GzLHjALt�/ �.�K�n����R�.�2���[WG���:�P�oHQQQ���1��̟���	h�,��|_��}b^Ml�5����CȤ�tt�;^��,�D=9!�P�CT�$n*L�lj���6@՜�k X�00X�#���j��xV2O���A�tq{��ـn��Mi����q��V?���b����_�!/�����wIo���h\���|�n�*޻�⬛�K��Ͳ�|�=�}u��.�'K������5�H�������Iks֭{�����I�j���-6'?�:�z,sȠD���
������GΌ��tF�LO�DH���/�z�%???,���b���dU��3=Ao.$��5�oX8"H;pzOd�Z�:Ma�g�0TdJkl��}��E�(��>Ǌt�J��S	ź<�*�Ű�����?'==����(BwGO�z׳�VL%xK��܌ML�T,8�-*?��`_��<�bⷍ�#k��Jl��,���<˧<��p	����.,�tv*�����Ơ���zk�.m9[%s�����Z�,��h�d..��3�׸���y
�=op:L� �����/�����t��^��+�=,ljj�zu�_e6&ig���%T7ZƱ���Y�"��߶P��6��!�B�x��29����s���rB��-&����n��n���ׇ�~�8Nx��֪PR�v&�啔�j���T'�~��mf�#x�%�#@�{s��?����
		�p�|c"Y�$�?ט9ɉ���[��c
����͙�3xx"�FIٌ�xx�)������r�B+���<#q^�*���?������#�bhci�`~{�h(1��e� a�m �
�.Zn�1���%}g�M�`�ndl�2,f�]�$���߇=Uq2�'u�jJC�rC̊g��D�����&���`�X�Nu�b����ȔU`ӵ;�n �	���ȓO���l���ڋ�=Y�̰P�x{�z����&;gWW�q���Í���\τ���Fi� �$Ň����'����	X(>�����j�@�ajYS�ov{q����\��֓���3DD�����f
�P��@����7ѥ477�U���J�c� �癹C� �d-�T�k<,�ϗ٬I~% `�Yz���@�ȱy��nҷV�4����y Fs�� Z��Ѧ��PȳIB*�'�P�|��:bL2"���$���~��(��˨�Go�.��C`��bgk�Bh�~�{��z� �C�^�1���OX���m����r�]u���8f��<y���k��嶤�Z@�)|N%jFH���SXdda�Ԓ/����;;%8��]��z�|a��*h���)]�0�̈́�m��ى�
�������F�bCR����|�в;� SS`[�Syu 8���F�G#��_xNY�����<E\]�I�z#$D�.Z=o���@�ŝ��ǪaR�
Cdh���[���B�[+b��sw����Ā����qh6{��
D�oh�: 9Uk@���[�~J�c[X��F��;+��R�+4a���?���ð>ב�D{��d�?:���f0%���1T?n 3�.�KU�dD�n2D�/on��� 9֜�FDD}����@D-����_��X�.%h��Z!���������G�f/?�{��'�]z���������Mqqߙ�mbu�������!ϳ
ǹ"/..�@�r>���6��;V���!��8�C+h�ȯ�Ȩ(�3�O��@\+t_^N�0[����Sj���ߝ#;9=����Y_@-��]�Q���:��t]�5��EĪ�j<�d�q>����]�L�8��+���2 �Ē��@ �2�:jj�ȸt�`0b�:����@h�/��e��(�r�C�	ڨi2#��B?��sU���Rx��O�W�;���i�Y��/�\`��=H_�9�R�wA�G
��Yt���a$\e��I�r4o���k�!N}��A��2e���@��z�&!a����\�M��F���*�#.N,�_����>��,=�����p��[=8��,p\T�>NjY�4_.�v�n���daH�?�MY� �=]N�(:Z߯��� Y���h� �bw8����[	��W���4����xW:�с7���H��!������w�+�a�����Bp�z@J�.4pN`c2�,�r�Z(}��V~xc�P{���ݦ�������t��N.�[�����<�6��7s�����
�8H;��|R�._�H��_���tr?X2�s��c���Z�4��W��,����z�H\��fʰQd�Io��ZN�/����_&�p��WQQ��QG|�T�g��pm[N[M�f<00 ��u>SiBuI����K�x�OT������Bm*b�̦���4�:44K�ru�]so"�~���i� d~7� 8�Qh�).��bJ�,�T�^�D��q_����o�C��{)��&���q�?Ť�)���i@%����X+533���.�˪�U��p��&	S
� ���xS�P(sYN����Tn*B���p���� q1�����|UT�мA��33� ��Q.�7�D���46ŝ� �4���5@��"B�� �	 �ށ�	�ޡ!z�<C��pgݮOr{�_�Z-4ġ4ZL��ʓ��� ���ֺ�4���0����1i��(<����q��Y�A���%��9r�js��/�hY�^������db Q���eC:Sa��_��!���ƭ,�OB"����
::���KR�zh�a���g+&��?��7N�W��zq|'zxZ~���o,cn����^9�'�j8S�]ߦ�s,��p��'[��4�y��9��On��AS�iKu6��3!�l���9NGI)�o�o����B�1V�����Z���f;%�m�G���D�T�j t��MZrrјP����Ύ$�E�����|���Nn�n8Ϗ�)���c�A(���<C>��c�Z�qĥ�p8�ݕ+Ѯ�������z�#[1���'J!�7J, #�bWn-�m�i�:�B��?�2ۧ��bP	X�V 5�`r����veA�pR�7+�����y_�P���آ��=LP=hM����0	��%����,���w;�ۃ����cK QB럌�ίw`
ź#�T+��8��;���q{}�kԟ?�L�ll�]N��g9%2�\�Q�-�"x���J3�\]�����\���j&��?���g�j���b�wGP�J{<Y�
�ٛ���#=���o� �Y{Nnn����Ϸ���i���y���Q��%�Ĥ��s��@~񥃔��0��8���<�l`��5n^���?�泘-���2^��>��ɺL�)�.C��Pz)�	0  �R�g��uӅ�h��p�"�pjVVVr�'~JƥG�2U�%�/�>qsq��"d���5���kkk��נ��z�UfԮ^'ɭ��=��������ӣ�~����V0^X`��@�gr��S�\=$�h˶���5�͜֋)@�v�I^�j��k�#�א �����?6	0Gb���K=q 0��C�9~��/���W�O��k������ .<�	�V1�yn�7�^�~m[a���vkdU��P�'mm"g���i�+++�D33$窔�&�����𶁹�TR�,�����ws(]w�/9�t'��v|N9�O�G���+�'�^���B��4�@q�$q�1ى����+��+3���k͟��C�B  ����4\�iD���j��+
Ί���`*|&���66�`���}�������	q���Vn��/<2i�%�u�tAYNc�uAۇx��7���ߔ�>��m�b�����F�ɐ���h��e>r����j���JW[��ȥ��Q�P���(���Q�l�E/�^�K䠵1iB^
��aL�w�|�|*T��F��L��)�)�g��\�~x�;�����+%\k�jӻS�1 ���b��<�s��U�n�w�r���K��#S�۾�'��m���XlO�sQQ}��.�X����m���ld{=>��3�����\�f+1��p�*�����
����<���JGGg�|��#��aw��&�uЉ��S���onn��Q҇�o�EQQ��lG��]�͚�%�����N�Zt��Co,��gJ0�^��;�m�ʖ��+���1�@s~�XX�^����C�ԙ��Y���R�'/�%$$���XDR�Rȧ��; A���`��.�}�kC����ӡ�W��4{{/|#��S���iҁ ]����p��ϰ?���l{�pg47뭪��Ϻ%Q�6�/}[��-�C�5����R��z��p�,��ݧ�-�/��f�/�P�_ e�k�����\�z���Xw�4 ��<�ԟ��Y���xa�{�d���5����+���{L���4đ��������q��4~&�iG1�M��kz���B5�����J6_jj���Dl{1轘�O�^�ے��; щ�bO��&逷��ƼAd���ϸ�.�g�$��_�J�grn;#w��X��^����Aʗ)����QV�����hn���+�u��B�����	��I+�Q��Fd�A@��3��7�S%�t:@$��Y�	0����s^o&[�O��3V�$ W�����eD�3g�&08���;z�����֖���~"�$D�Aƭ�NWH�䅃�|�ԕ��dal����?��+����Ȱ^lJD���� ԰�w|���7���(�@����t��K\�s���:"(>>�g�b��l��,	ԘՇ-�����`T����ҟ�6��������x3W�7�#-�C7���Cyi/���+����M)�#�C�������$_��*(`T7������ja��Wl*X��}�"�Њn��h���W��Ł�f������J���۟�d�VA�nO�R����H�s��c������~�����u�3-�'حvp�+�Thli���`�E��ҧ�hs'v���y�kEnrrrP�Жl��2���;�}ꌬ�]�RG����44Ϟ"��r�߬X���;�k���Sw(���2��\	���C���O
��]�Ɋ�ͪ8hVw�

�_��i�t��J'�aD���@�&W8�e�����^�].yIm�_�Y˕��bc�@���� �d�V��������`x��_��S��k�k�H��m}���LL��f�zy��Xߝ���]�{��s_��?�ۮ�N�*�(("���DBA���-17��z��`9��4Yy{@���tt��B��H Kv�|_���W,�L�ٕ|�m'qp*C5_����ŌMF�9�2�=�in�D��Ƃ�t�`�򑋋���f$PW�~����x���xaL��O�5��F'L�����EH��5������Myh
Ϛ�{ �#?oD�e� P>o���ȻǼ�C��!�鵇��{�����;����{��B��eK�k���A�޲g��*�-eoٮkvmQB\.�k�Ȋk������T����y�s�u��9�y���>翯5��]GE�j�Ꙭ�T���M�B���Gl� '�G'
~Z_�/
"ᖇݵ�60z4{�!0�)��sס{ ��8������.����9(x/���a����� �|38x�/��Cu��������YE�BW�EB�D�v�@@R2՞xQ�W�����,!��*�:000]�k�*aOq�]�=���
��TY�`��-LKc���*7aiShp01p��1����8���@�"��b�����==�%
������A::qެ���9�U늇�	W�	�Q��]ZT�����F��0Z6k�--v'��4=3z�{J����q�Ak]���k!�ׁ� "!��M.I_�x��x����+��6-5`@f��D������cN��OLN^�ї%w]S�AZFF�2�<Xx�A���O���'O�g����������=���C>���~�g[�X�N��A���	�z�Zv�5������_g�q2�B�Ѐ��}oo;�خ�ޒ�0�����^�)�9olx���������	)��N2�������޶�=�"2����}���OCF#�G��T�W¿#A���n�����U�Ԑ����G'^f`q�C]w�X����ۄx��2�Ɨ �p�	p��k�	�\!��cwѢ��W���}�,Jl�%�!�I�IH��ߟ����~��QQq�9��_�$D�����Z|��C��ҨB���)'�i�N݈Rhd�_X(p3�����Բ��J����;w���$j��_��x�˰�<����`iP>F#�穠 e``�+Sr�\�4U�����*7��c�R�aǲSs*lFk���f�]���e��UH��i���o��;����^��h��ŌS���w4�����U ���mAf�����廐d���V��'��o���!7͆O�E<�ǳ���FC���K�>�H~���P#�՟K��������P�MR11��,�TU���g�%{��;'���w\��q�$�#��ϡ�Z�s����A��C�<��!�M�����?��NT�yM'�j�_+�H.�+~���kԕ����5Y�n�A�_��Rr~T6���݆.�����o��\�2C��[}3�J�s��߿Ia�����&��c1W�Wi�<2���`F�S3�N������d�L<޳h(1����俑#X�b-���;����..."? w��BJз`���}u���*�N�b|z����9��� V�>@��43sfqE���i'`3=4�&Su�e�W+[ۧ���j�~�`�Jާd�k����T�sVFf�b���hfm�Y�tJJ
��*{����K���k��.,����.`�	!��J���{̬��e;�$�VT�sנK���q�b����׻�ty۾D��F�E�a�2{�ɻ`B�����O_}�ޮ
V/��Ą��2;(W��������]qTU�'�LE��N���V�%p
��qʾz���^��O	��U-�ͅ�/^6�7:�1��mu����e�P=3���6��[���N��YJ
o#.(��Ǐ\�Pʪq�~~*�9|�*$����~�B�Of�P"����=�H��`7	�߾��	}�]�Z�f��&g�s�����_z�Z399y��)����9�R�V��l�9�[EF�U�R����ssq��|�N��|,�h�e�/�p���z�*�d{;�TQ�joeO�W��$l��P�&�@/���gfƼ{�$x0�ry��/<��04�9:9�ZK=��a���mW�F�J�~�MJ�2��@�FG�)YAAav[������G��gj��4�s���̘�6�|�"���EG�Q�]��8\4��A��/�x࿭�����s�#���Qc�(�QM�'��Z[�����1������,hv�	���K��x�s����w����A�P0�T�0zll��,i�_�	D�˧̋�%Zq�"�����퇧�9	�*�
dKt�c:�Y�{��nnq��W�M\]/�gdXWwEn�m3������>'�.����Fz~z�8�h��#�1Xw��ݚ����g�(����R�"t��	&�/�>���9�����l��b��~8/�s�a�F���`����[��c|�Lt,"
	��bZ���٩�8zB�=G�5��w	9G���4;���M��`n��a"������f�d�:z{i����lI(���Z�qXDB���$��S�*��|d95o���8<�$|�X�Ei0e�	O�ហ�CB������@�Q��P��e�5�M�N�,���Z�[�˕F���(�]y-��&�F&�<5(l�I�BZJ󜂅�d�=��/��������X�E��X�N��P�w�~��J���@?0.��� ��8~TjR�524Lߊ/�T�Nޟ��6��\je8�@޶�;����@�`�h�b!o�1�#l�� �/�w�����NTN�*�]�7���B�������W�9�:�+8w���#�P�Sn@��/�w�0�c5�8�J�J�������W�7�g�W[|��7���t��c~�wUv�ڏ��?�w�؇�8j�o��p����-FA��J�f����b|��/���|\�O���@�? �W��m���e^�_�@�;�b�G���'ֱݦ���0G7u�vTZ�a,U��`�.D3�c;������~�HG�ev�Il�D�l��
����0�w�%p2}�ۭ���2/J����$�nzDfi�F��y�z�<��ۥ$��E�݄���CЀ��˾n��3_�p�Wn�o�����t�/�������gb&J�WS�W��򒘁V��pV� 	f�W���/�0K�P�"SX����MDx )\L���kf�o���S����Y:42�ݼ$q�Zp �[<��z��J�{bQzh����)�X�*�����qӜ���d����Ғ���e�!����9��L'�Q�b��5Q�ȱ/����L2��A���:��?_��?>Lg����S2�������=~���t����� N�����#���.����� yi�N��I��>ۤzGM�5w�,7��II����O�>B�D�K-S�j��*QwF�,��@r���ם[���o�~�!�I^ggg��W- td|�m|�UHH��������G�G�)��g$$��_�}1�L�W��֙�E�A��Z^ �	���ٍ�$�C	0Z(�Ũ���kB�nl�����&J'666��×*�_�>!����-]\b�P�R���E�2���^Cv#�����MN368�xJ�<���"��U��n!Ϙ�OU3��	"\?p��h��E�m"~���j�<T�7Ď�%�����2Ggf��vR��iO��dY���Ѱ��P�uj����}��F�S��=C]1��d[	���3-Q��jC.��yg��=�;x֋����拂��0��^(ҽ)�5�������>qRb����������3WlU�@�.Ňߧ£!a�b+sC��9����Ӊ
�;��k]��I�+S��<���*��K�S.?�r�!�++0g͑���(�}�9�	*H�@��$��&D�E��
գ0{L]S��	�EfP<���-(�@�'C!{あZ"n/�lF3����IW��y��:���}���]��*�x�j&�o�1g��|=��%����n�(��*>�0�OJ��XMZ��U�OyXօ�+ޟǜ}K֌�R���ܸ��,�r����ڿ"?�z����6k����@��Ch=�A��C���^0g�C���?���V':���fF��$#W\]C������8_ђT2�Z�f����W���/�)�K���񩸰��w��^!-���~�rb\��Oʻ����̫�N��;��ك��:��B��K]YhuK?Z�/_��Eگx��-h������.�r���;��
���K��I��\���7s$�D#O�,�yW(1�$�-ż��c�f�p4��ᕿIl�'om;Gd�T!������#�+�	2Z�60Lrp��C���
��s�	�gP'F=Lc^�uXx�gf[V}�
_�I}�,>G�+5�"t�7�F���k�@� ���M�.֏�ȓQ���.�³M9����y�ٺ��ɂ �(��K��3��}<�|e�L�d�1&��/�T"�z��8��@����u�r n���4���'X�`�7T��VP�����GȒH�S W&��m��Q�w��I�A��6os7~����C͐@�:��~
.^GWr�S�%�4�๺�l�Μ�o�d�����5�"B��F�y�~o�C~�jF�9m�6�3sN��^�Z�Dܽ|5�4:1�%(��st�,7�|@Bo�)�R��a)*� !b
1ue�}�h�`�h���#��ʡ	j9HQt��bܦ����;;&I�3�VGP#���nT4�8�+30r�,�!"y,���0���8��85���JTq�Z�������K?j
2��#����N����:���e6:��܋�����ou�l�3;e<��8y-����,�;�Nz;aZ~�g; =Z5q
�M*a/ )�4��2������x8���N��)��\ﮩ@���5�$<�n-������L۸Z4u֤/Z+(����u�b�|�}�|-%�m��V���#!�t�t�im�}���x8e24 �L.u�Id�\+�2���
3�OdA��rZj�M�֢y�~t>0��T	�FQԢ���ٽ��B��n_z(��P��v׉���y�b��3H�T3QG�Nvp�w{�Y���Py��͙�b�����0��m>����epҠH�˵��GrЎF��Æ��TfٰA�!/#����5-q�lQ����K,��R(O��G��|�V���[VFe��Mh���,c3����"Ϲ3��j�O��)bW�e����.�j��!C&<���f}G;����}�@���F�ԱL��@{����e���Zv�1]4�=ތõ�6;2lY����FY����;k���[j��A�A.��6n,hO
k�X��[I��+ق��6�[�5-<=0��C|H�7���ҹ0��&0Թ����H��������쯺���G�K�,<=?�oB�(�M�s�[�q�S���8^�L6z��>]%&;H39�ٺ&�͗��á.{!=%{߿CmV�
�ю�_B�G�L���{���������,]]�ǾM�e:��ƣ����̭Q�5���k�>>#cߞ�#-*UM�&#���[T�rppH���=s{��F
�A]�K�K�Z�!CO���<����w�ik���H���3�m���k�nʋW#�����aoO�K�K��V9��L���YS�c$vA_�}��H׎�S��F�����?:zc�� S���E��k��_l̏��.d��J*u��r���N�����M��ݓy�����x���V�_Ȟ��?���5��[=���5Ԭ��,¿L���>y�e�!�����R�/�M��v�����<�����-��͛�Wi׾�άsŲ���[�
�-�~R�2(�3�8.{?�}���o�_�-����=ſz�1���n���"k�J���`h�����6�Ot�q���a�>�@+I=^���Y}��1�L+��������J�w.�IZ
7=Q�+�kh�hl֭)l��@1�FGGW��X8�f�U2Oe���4)-/�����е�'
0t�/����yR
���h8�SY2=#%���BSWO����C��J�����x�&f攌��I��f>'�MuOO����v�n�Ӽ{���� S�fqH����/z0��6m&	5@q[�����Ɓ�SQQ���=l>�TU�vuU %�eQ�2���q?Iؔ�-@-����.��326����X��;II���#ͱS��y�=�P����hchj�8Q�a�7SO�wہ}G5�i��ΘB�).~g[.ֲw(��MT�::�mmmY]f!������G薻�j�����a�K���,~����w���X���Q3|"�r
���->9�u�Ew	0z<L�F���hUq������h�^Z�T_��#��鎬
g�\W�d��kq�;f"��h8�2� ������
���G��{�s���)���G=ۇ�Ѫ��e^g�V�"����MC�6\tN�l��+>Y��r�~,|�����Բn����S�m�S�<ڣ���3|�]�'˼��O�G��@#����)o㤾E��\�H<��Ul����B�.���8���@�����\�ZڦR�A�MKN~� �Q,Q�٤F��~x�~r9ڋ�����ى����s{��+d04Y��&鬯���0����e�5�v������{;G���M����y���B�];�w�f�V�\��$%�c�@��_g`�qtq�拾�*��H=�Uڻ�闣g'\e�F%����
�0���s�a�k�;£����'+qS=��������St�������Ɠs��Ϩ�����^4;iC��ڌ��հ͐̼� �&�lsB�b�Y�Z��Q��:`(�1������f��i�m����h�΂�/R����)�tV��{�@S�e����j?��>��ǙG�٨ �o�\E�DB��-�������`���# T��B�e����lΐ$dl��r3�XS���y�0ws�������2N-_�\� (�Ru���H�~��|�y���ɼh����R�:Ph&aZ�����b�Jۺ��H`T�y����.WA��3 m8�����Y�L\]��~Q-���ⓛqS��_���C]0d �(�5;�gb��6��	[���F��5�J�f���$O�<Y�A9q�#y��1TqS�`���I@ R��fXT��xGn4�q_��L�m�6x'\㠻����0�ge�$�CU]�C���Q��{����=v�.o\�9&�@�}�?��5�ߩo�>IV��,gt���#�L���Kg5W�ӻ9�0.+�
�z؟ܞ� �2�q�T��}�l� P&
fv�� 8ݡ-
��Gu]��d<+}	݊h�C�)h�{�$h�@�(`4M�{D��r[Z�l3}�=zE�/K]Wx�+�����������cb�2	j�j��P��1l�{ͱ����'(J~�I�ԔsppB��Gr�+E�X�����
~yT�Ogf�׷߾U��z+����ܾ������;�^t�0,�vp�(v����Z�0�x<	�"�v�tWε�0���9������7+���b^@żT���ɻ6�Ȭ�>�ey���>B��žmz>L��Q�/�b����c<���
,��i�.�$�66.������p"���Z|ʕz��0���

��g��.�V�:ۄ���<��j���w[�w?���;3s���/��]���d7���՘�Enk�{��e*��B�E�ylum?�iGk+�3����v���{=[�w?L<^S]]]o���Au]�}\�ԧ��p|QB�������^���{EB���y�C�W�XJsx8���Ji�1���T��R?WGG����~59>�?q�p�a�f4��ȥ1ћ��el���+sss�bcYu$3l�x7��f��m�������;.�.���H����R�NG�6Fj�$�������[x�m�>��H�|�p���t+W�K�	j��CP���nWE�-�|�. ^�����N�3צ�or�=��LӜ��Y��+E�z^�V��z��6tgw!�W������J� �4�9at�>ށfP�(F䤅�	�WY�H��}n9L��LCO/��5��(}�%C:��g��8������1�*g��M���<$s�-Q!,7�o+�)�=�PK   {c�X��g  n  /   images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.png�xUP�u��{�;�)�AZ����C�I)�-����8��P��+�{���tw��Μ93�pfv�,B��*�  ԠJ��&��q��un���j�	 0�����z�Hj/�w^z��^�V6 ___>GOk+7>W��S) ��AMI^�/�$���Ġu����������1�6�b���w ����(:��9�A�B`hz/�抉���T�K����%U�0�2!54����+|������#�lI�)���ŶE��V�c����m+�h�@.�����9UF�*o�@��Qt&��t�t�DA:2�L��K�H�e0�j8"0��h�����A�a��/�b�V�D�o��휞�H���l	}� }L�~���>��t����|f?�Y�����0)�){��`��o5����1�䩩��-��&�{�6�P��54v�J*c�?Ν/�yޣ���;_�����WF��� �z����ܻ���1)�?�n��9[��j��U�Ҫ|[;9�K:�D"�m�R����7 쟟[�ެ�68��<Sic�"�lM��ljn6b:m�&L��}�pj�������\����ֶJ�U5�tޢL���n�l�)�ox;nx�TY �J��y�I�@��y?E�ʯ���zZ�Ҍ�w�;��T)�?'Q�63�������W��:�@��e���4�R�I`��V��ʿ׋[��^��FS��'kc��������k����$C��7HY�T���H�"n���v+k)6���2�& �gg���;�>=�y������SAJP��f,����ׯZ�:஀[�?�q���Ǚ�UGtY
~s��^�F)O�\��Ý.�`{��3��b�$�[��H�:/7(���D��Y4�zV����;�r�w�Jtw��t��iYuI��>~ɺ��%�^4%����o}�͊��!b���k����PP�N�˺���y^�i���	?	�<��횇
���<疗9ϺN�s���Y�S�nF��r4J[���松>���]!faU����3�:ːG�q_�
���?�君���g��fٮ��v*�	���P�������)��Wic1�&��
�*�QB�#}�,���Jt��Ut6�c�Y�RY����m7�dgF����w�9f`z~���������4�)�n2~��m������遡`W���g'�x���!���+�y��Dx���/ǚ솎q��0�ط��S�<�+�/@� J��,jnn6�FB�YW�1�z���0i��,[����zUiQ;�D���ϽL���HN[��|o�����\m���UU����@�Q�������g�3Y@�/���Xޏ�w;�s�n�%߷�WtMfI�0�c�IUr�{��K�����a�u:S�a�n|�IY��ARĈՈ�:� ����;4�JMP�64���g �6\]a~��u��E��5M�e)����N;�Y���@̬�{V��ɫd}<,�� rp��!wL]ה��V��`�|��L&�E��LJSKy� ��V�;/�w#����(�.��o�L*��P�,���L��f���n*��/f����k�M��C�I��V�{��f�9��e��x�Wڜ{A���S�z�}������:L��3�DR���5s���l��x9�o!�b��9�!��9�����ӖJ#v�2w48SݷwӤ�Y��VL�kR��NX�I��w�L��/�����}��ͧ���^��hx��x��|Ԗ�+�鳵�	��H|:Cu��*Z��j?|8c�{�|N�1)���.LCCSu����L���(���(]�:��@-�/!�7�?�X��M�-�p�.Jjߺ$�s/ls͂��Eg��L�8�:�?���{t	)�|��V�~ܟ�����n��Lu	�gAOB�����Դ��>
�g���xԂ屙�WȖ ��#�!��{�8ğ]�7�F�G}^���8�xڎV+/��f�}�X��}�,�<cj{h,j���~f��gi��Z�陟�`�c@�3��8���`̂܇�7�7+R)wQ6����"z���:�*��F��7�|l���nI�o;u	%�_�ۛ�?>܃�Ѩ&~�	 ��:#K��6
n�F���4epftg��(���Қe��M�o�#�a��%�:$�O(���SH\'dn��DN�O�)�Y��"<����?c�Ǫ���	Y��;���ª;�lH(�)x[t"�"G��<��㬖�r®�k0�&�`��C.�"0��<e���a��@�^�c��",N<�s�9q x���f�\WOL�F����j�&l�f� �����0����=�����	�@L�6Y�Ed��Cy]���N��5?'?_���Y�q|N!u�ʜ�s��u�N`}���$~��g��^�z�qr	J^b�e�T���ouVT6 R �zynZ�e���ۅ(�0���ȗ�<Y�/�hm�K6`ϓ'�L4a4��{�щO����������"�M��8�;>������m+2/�O������2xS_:x���S���P��A$�޳�l�ϞY�(���5��l���M�'ק*������w�}�����Zq(㪯��ϣ�,�݄1��-����E�w�>�k�O��$ܗC�@x�j�]��O��'N�TY���"\���Q��K�iJ�y��1��欎|��q��b�ӽ�#W��T�Q��ݪ�6�E�#g}v�\|)&�Π��!��S�y���k��i�$��f�*����˫"T]P2 Ȧ��$-t8�j�QG �7��XV��#�{��L�v�&g|�|�;I�Q+>T�f�b�+��s.�	�]t�ۃ�cm]N�û8��z���׈0=XX���8l����=�]��x9��^$9�m��r��/���Ɗ(Nwn��X���Ea��z/�ejǫy&�G�A�1��u^�U���e�Rv��	A���L$��t���k󴊧b`�x�`�`m�c�[m|�q����%�`���tl&i��{CwC�W���v��3zB��/�0
�}���j�FχY�e��QeUNh/�e�违:����y��',�[`�Є���l�#�w�-ܳ�ע�yRx�DE�����.B��l<զ�	�b(Ι�O���5i�K��Վ���R�'C�2��Ut��v���R-�U���H��Sh��W�\h�a3Kf"!N�PyMlOB��	��ɦ��T~��p����&��.��`�|S�����YP�H9B��7���'67���!�2RT��l�K>P�����F۞)/���� y�I���I� ݺ�
혷7������v���4��YH��V~8�(�y�E�l#� ߄ϲ�̲�'7@�eV�M �:P�����D���U9&��*(h���p��`�V������Z��ڎ@����Wu���T�xhT� � �ɣ����w|��n�X����7��`���PI�l�� ���}�wd��.�Dj�z�P�1�sB���E�!w���Q�(�����z�Y���H��-S+����D�Gb1N;h	���4A���	��73o��Z/	[)*�PV�"6ӱ1S�$RϠV�+��_��A�>��2;DU�l��
r'F����m��;d�7V�+�YW�H����4��5K�/���z:©��/ؐ�O��n�w���f�eD��<}�?�Ҽ��_)��dz����"��Y(v�+cZ%,�`�UH��(4���ٯ�P�e�+�靑A*&�4Xf�%�#��#�(�C Tq�j�YSu*r.������K�<>5W179>G��gf^~�Xݹ��������.+Ը�.��� �	Y&Ic0mu�]��;LlV���ֆ]2a.�|�K�FE[o=�a4�X85�=�%�P����V/AK�Ndb$���
���(2�R��t�b������ޜ��R�~�kbs�ۦ�]�{��&S��Rk\B\c��#��o��x��cK�\ۖ�1̥܊ou��p�rZȠ�xu	焝��9ȟާ�F��|nG|Wo�bhp�Y��`��sb+����IK�h�=�6{Ǚ:_���������ߍ����B�"@sMGK:�`P�Q��Ls��A,p|��{'�ڤW�/D?EWp�c��؊�o9M��
��M�'�c�{y�z��e�#�F�l<�B��]O��%۰O%��<r�e5C�f_��!>�ν���g��_��/gL��f�#�EgN()-#\$�\�Y���DB>'d�f��d?���@4�7h�
ǉ9���x�5�������:V19q���WxQ $���%��56��	�2��ea$�E����Ғ	�tlRh��`	d-f�Ԓu���:&�h�S�3��я.˨��v�ٜ���j$cT��	�$7~U4��Βy���&��=���Y��!1b({�o��rz3Pǌ�:֦�<G4�R<E�e�̼螪oJ�e�=��{�ތG���#��Mx}I�����G���1[g���X��p��ѥ,ߋu�e�&N��<.Y�WNH�k�|c?��M�
�t>�,�s|�2#b��-j)�������o?�ǘ�}�U�ˉ�V.f^��q�`x�9��K�!m'�������7�-�QMs�E�`λ�_Nz3
?�;�e�͊��~�]T$r�Ɗ/U��
}B^���c�k���~���7�jF�.l�g��^pr�3��+q#��)������{�{�H��C���c�L鈈�B��\�c���ġ��q���jh���@d^�Ѯii{���;p��e}w9��l�����YT�'_!ߚ;���¥HfH�+�2k�5�ASF�j�ʙ·P:{���s��	��d	��pT��!i����x~p󂭡�RS�R\o�"V�XLq/	@�U`,0�������""����*܍u�P�xC�|A7K�e#,�b�m��:��*�8�NB�������X��[���J汁w?���h��09qװ��~�g�(�5�׭�F�J���_�J���b��5Ƹr����z:P^��kϹI��\��7��������%��|�SB�/�[Q��"��ƚrK��T��(�R��T#����-K3uwUi�4_I®g����x��t�S$/�������v�"'V��c���)ʮl�R�Fp�I�xrQ'f$��[������X�%Z)	��t7^�RƄ��g��:_�ޘ�K��������.���*�|�!���K��s�?��Rl9g����fr��F���f��J�CrVZ��_�S���!�Q�̛��D'~�A����W�E�pP!.QC~:�/�y��$�c��3��4��֋��ULM��W0Q�v#�C/�B�9��q�=�݄	 S���E���}�AX��a��*� WMa��ə�qOu���EDO��k�ء��NF"|V1r�>�R�ʨ+1�T��@	'��x-x��ˏ�g�ea�{&z��6=O5���p1c���X+���cQ9bǆ�����dj���[���d-*b|Hvցޫ��i�zeG	{i�*.�P�a*`��!���]}߷NM:V�hR��~�
�v$|�RP����(����'�c{!��8�[z��!p`�����B��۟�֚�-T7!��0 ���A�Ԑ��@�$�9	��#��AV��ZO�TL�����N���V��@�2�x�M`�w����@T�'��B|�T��)��J��o��))��9)ӢD��s�a�!8t��le�%?'B��p���?�F씿��������_6_=UbkN��Mj��Y�d�_|�{1D99k6��Z8AM��ƪ�����rF�Aq�� MWZ��m'FM����;-��<|��t�mN��a��O߰�O����O�',���;_�h��u���sm��$W�S�HĊ��ԅsv�wث
�� ��2E��4���a��y��ܖ���䒺���x���X�>/�X������w;Q��kG��J�ի�q �6ǰ=��I�u��F$���س]8���3�F�j��)�/!ݲr��Ք��4��l��hgf����c�&�IK��6�!�Q0���x=��]=���,��d� ������0;����=��i�@w����sk).�sOvA�y��W��oh��6#��Mbۍ	Fm�����F�F�2��PK   {c�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   {c�X����	  P  /   images/471995ad-a105-47c5-9945-45370623043a.png�VWTeai�R���	EE��Pŀ@��P jiF�J�J@�MjB��B@:����Ĉ˜=���7g?������y���n*"���17����!X����t�qfN!||
���/o|�l��xcG�-�O@����o�_�'����X >>�ys��]X�z�-9�lI޴k��5��v�T����L�T�>{V��6���褠��.��cG����aP�]B���8(M�L0��s���@�Bݔ.�tQ��po�W��_����A��ނ<�5.oxW�1T �ӸӮ������Vi_=� �8G%����4�"�c��(�E��^G����"[�#"���K{�k�֧W��#&CUr�E�����޽�X������\�R�8�<ui��m���g?yg�N��[�4I�g�766V���w�I4ՓB�"ٴ�ȭR��(7ooo/U�����H}m�FM]�jE]�<EEZ�-ӳ?żg,��!�@�̕��e�8���brI�^��|.���Gs�j�Zε�ow�����0�l:�l�cCB�^��\i��}YZ*��.��dlBoRj�)�L��_$��{츑I@.QC�b���>�1��ũ��{B'��'�n�|�����+=�v��U�60�M�y0�M�Y0�4u+xa��T��U���>��<����	�4vw=]|���%պ�;����}����o�em{�J�Vab4�����F%�f�Ɏt82�i�e@ �P���Eʐ��l��������èV�M���\c��$uI���?�;����˗��+�se��Y� (�� ��e��<vr�/#����۬h�Dǿ��4�z�Yx�Kr�'`���z.�Xb��4�\&8����?�g�^��j�*��@'��%��l �����r?�}��[p>���_5���2^9�G�VQ?Ӗ�� ���:_��?���eoՅ>$��gըOe�	H3q��9��G�?�E\B.%�m���D��K����r��k����e-�b���)���m]�Jǩ;C���ӘM[>�o��[�Yq��#m��ʏ�B�G��>v�gB5��?i��&<���������R��G(���l�eU��i�$�����Ɣ�|�W��H�c]�Y�^ubU�6C�eٌ��������Gs1Vަ)��e�`_(t���"n}�����@�;Z{*�C"���P���v��H��sC��E�R�����q�5��ee
`���^��j��C0���H�́���_�{:������i �ɱZ�}�ibZ/�3!-���b�n�!K=�V����I�h���BG�#@����	?֒���Vl���t��-3[�?�.z;�[1ѽ&��]t��J�_�7 '�&��}�X���;2%�|�D�ӭm�;y��U�<{�+T^ZW��A�]<�剠�B����dxs�5���I�J+�#�u�>��]�^NoeM�^c��(�(�2���a���{'M/���{�ɚ�$�KN���5�W���v_|NH����ZV�,����\���0�(jA*©�)���8 �1�~R��j�����x�P���{#Vm�>@�\q�Z�\�mU��N�~
t���c�VL�������q�a�9��4Sn��`%�% )���]H��Ly������	>e��G�O�/DҤDL����7�}E*�l7�t6=�uJ=pO΢U�(Ɩ;�@tsM&ہK훬wOU�y;����f�%������k\���	 O�n6dBth���3�Q֜�+��#�� ��A:�~�~A�<u�
'�R�(�i7s4���VM�$��;��݌�;ȭ/������ȩ�"�
��b�w-l��In=jՌ侉ڡ��ED��G{,�-��O�ɻ�0�l���%�˗c��+׵ًm�Q{A�5B����u5�ͧg$�#���j��!b�?6Kq���J��3т�����m�8�<"���>��N��$��d߶�;��7$"N����;]x�It��\c�Q����m��h�z_�f����2�:��ԍ夰�����عH���U�m���h��V���W�����������&t�,�=C[y��^�$!2���������u��EVs����ᮘp�Qղ� (c���U��7a��*�����'����{9�h+��n�x�ۈ_������əwg̿���(���9��?�V�L�$���A�w/��Ƕ���~IN�?Q�?}��[K�����ދ�Ĥ�Y��lg�
�� ǂC|#c05����:ͫ�Ɲ��_�%8Y��Jyv��%�-n����j�e��ؘ��S�!M}^�N�j?�G��Uj���}l���XOZ;�;g_�FL��Y�-0s�#�[��Θu�<"�wv�f�
|BS�wy.l�[g �l�/������VM��iU��ٍ�m~��?]����׋�gn��A���PK   {c�XhT���� ċ /   images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.png�|y\����Td�D�+!*ZD˴qk�J*E�B(�F��-��"d�V�j�s�!5hE�(��}�]gD��<�>�_�^��m���s��z_��u�3~�5�7od߈�`6��(��`60ƪ���/�싿��8����������7ت�s�`v�F��)�����vCQ�������/a��Z[:�_��$dcoE�a�`x0�
�u��}�R�8��w��`��&���`>�kq���x�i����-�S���q�A�rg1#u�]�u�\��ʖqѽ��D���A��뗬M�N�Wj��S�1N�0�����^a0-ⷥ�^2�;R���@�z����f����n��=S�u��x^����:v�5��+�5����;����w������;����w������< �M����R�̼��CwR_y��ح�|2��t���S���]o�[��}��C&-�Y�5�	Y|�F/	}<W�|i^u��b�ud�MK�e��W1�F�]����F�I�G������&Zꅽ��c������7����Ϳo�}����������lY���и�vKr������?���dfE-���aƪǛX�nd��z��"��&�99����]�ʎ>��4��u�8�O �d�%���	g�}��&U���x]a��{+�;;�٧xՏ������ZB�����A�ca投�B��䠏����d�������l�i
^�QHȤ�����[W����9�9�nj賍q����#I�_��Y�6l���xrR��Ӯݙ���\�/_�Ħ�:�|lB¾���FB�q%%r��~ۄ5�*����i;�)B���q`�~�*���;gF��:+�l<�'�%o�9�I�?�w$�+j)��˫�,ѺU;�_�vRU8������Z̕�~�!rMG bf(��ْen7�����^ &F��}��l���^
�ŚU����M����{���M�yWVRPPP2�9A-�s�[���4<��ʕ[����!ܚ�v�������lb��ˊ������x��e���fii�����C�{����ޘ�׷�u}xv�n��Z�iĔS���߄{ƣ��yL�Q�'L�9���\-q|���M�99G'�~�)��璛����Y6%-y�c0+� 6&C��uO��\v�zK�W��a���[k�L_���g����sRv��Ǒ<St�fF��d[h�J�l߯}Jv�OP^+5+KԺh�J�`{�����ʬh�}{��٤]&��oү[gnjʣ#�w�f(A�N��ŕe��>298##\Q�jtS}���$Q���7�|���	N�f���k�:9===���h<��uA"������o�aDј��\Y�v�
�U]�*�SSSsbb�≔C�An�U���vRڑ��k^�7ݺ�3���k:�H�WllB�ڔ�>8xnۏ?�{W���o߯Q1?\�=\<m�6���˽������^ϫݧf�^�L��@vp�4��p1���5�u%�m�B���뿼��/-�K۽����I1��$�]��WX�֐�J@���Z�;hTp+-�M\կ��r��Ü������~]�!I��0?��f���󱣃;��ACC,��������l��Us}ͳ	Q�J��`�mk�������\gF!�?77��au��[�I���%6��76oN�.?��֢e������b-��3��&'�sJ��{��p��;v�����R!ս����r�#̓㐣sRY!«
Φd����hur�����|r1�;�l���M�Qd:*��D"���rdY6g �&���^C6dQԪ�U0�h�i/�^
��]Anb�.��������?y�ĉ��Ϧ��Q��[��;^��\�Ӟ�,��_;:ǉ�w���>>"!Q�.B�+ڕ엘�H=қ�w6�t�,/X�	�}s����6Zǌw�ڔ/,--=OM�c���-����A���I�'z֐x�;�\&�KܜQ@R�.FL�Fʝ'�͇ۋ����b:R��Mi�;��)��L�� k���;'�MB��m������[@~�	FٽV�S1��Y��,�3���-	�'��j�Gf��ή��Q����RT`	l	�^�4�$i�]e@j/��~^��QQ�)�vLJFFF|I��.y~W�Ǹ��{�e��i�������335�M$J���6:]�,�4YZ�H���¿�n�E��SR���eV����T.f�}v�0�ݺ:C6��G!�Ĵn��p���Q%���uuuN��������/�Mca5�=}��o�G��~+!d7$��#��H��n��F(W��8l�d��G�V�8���.���˺֘�4����ݺZk:������Հ�q!r�,�"0����l����D����|�9MG�A_i���Q3Z�ɄP��������y=���7��[����㲑� ����Ӆ���c����m�/]�v��{�.��hW!H�g������O��:�8C�jr[a�XwM���=Z��;�vG�ef
���h�! F��-�a�� ���d5��0�!�sww�Y��ʺZ�x ��T�|-��KJJ[j/�.��h#��N8��JTfm�y�?��s�OԌ�%x6�Q�jn�'.[�TI�	�]o������ͩ'x/rߏA�-��6O�=�&�z�x��8_p����C;�ߣ��E�/���Us9V�ºH�o'��ЭoM}C��2�
m1Qd�c�b }��~�ª �	��'���-+>�����d#C[�j5)b�ޅ���e���G���V�E����mQ���7l狧v
��g�v?2b/�Ĺ�G&k�l�ׯݔ��dIOv(2!��jf����
�Ľ��h G_J��?��@ �h�Y�?�m��I�^[�{`|]�I1�ʻ��1�N^^Z���|���@E%%Y��j�^}��`q�����J �@��]8���fn�;N�'����������v��ф���1�@pnR"�6���O����z�Z	��<f��8���=�x#/���?~Fޑ�����8���f]�۠����SQ�v
s:��%E�%���tF�.\:���I��/�Ja���;[=r$ܥ��n[���n3ʱj�/�hhnN���Ɯ����oC!*~��A.��LG�[	h子2�����Q�uj1@F�!C�=���|�ܻ�.��5Y��\Z�c%�@o�:<\���	kD�<�/��ikk}'���o�!�v��% !��@)t@L`C���\��L�V~�X<�;�
V-�z�Ȇ[C.�?��4�Q��o4�p���-�Y�	6�cC3�V��M��� E��{ ��P���-¿��=�6�"�M4d-t�L,���jB��R����D�����Y�(	������$yp��+3=�<;�Oe����8�v�����Y��Gk7�!7�m�w��i6��D퀁/@�!��K�[�mpHyP��E�i��B����E�#�Kz'�nr��>���W7�?�]� >�������˓���F�f�LZڃRG��<W�~j���
2���]&�I\��^����E�x�g_L<�O����kF���k�a��?�4�z�y[��&�?��9ui��p�%'����uA;:Zͭ)K��Ϸ��C���X���NX>�P�D�:�bt�����#�~Jv�%�4�S �� �.r��^��B*��S?��!V&�|����(����2�b���kq��%�s����^q���T*?#jjj
t��O,�fVL3)�����F#��#�)�Q �Iѡ;��#a1{a�%b����J�|��q'���>���H	���Z�!R-[)_ʡG�e�����[�kܧ�X �թ-ɺ2�V��`������'e��i���=��c��f(��E(�W��sW=IZ��!x��g3�|��}^X(A϶�q����Uabj�*�(����4P��w������~Ϟ=kpeWt�?2ӭԮ��{��E��Ln�e��uD죭�(����KT�3����^:S)l�99)� �A�-�{��Π��?�í�կ��?~���Η=���CP��_�����"kFA|(��˿����dXN���m@��|j&��ʦt�8v�����r���&�?�OZ���lqn2�"��qf��r��n��v9��r�{F����wC��� F?*s'DN�z���H��_�����2L ��-RE�D ��m�	��8Pg�� �S�-�4�M�_�۾�
�7P�?V�p`rrr����"B�K��e� ��T�eg*#����l)�YR ƾ-h���U��c��xO�����uR	�8�|�KlT*�\�Fi�A,#U��@|"%&n�rυ�j�.�Ifs���qB�6��X��vC��#�X�n޼y��M�
���7W>���[%�l``@͘=fɣ�ň
Z��IW�l=A?v=0�V��?S�ɉ�
J��|TR'y��U4�jSG�JgV��ԹM�ʊ��/_��2����pE���p˳�ޮZ̈���{��1)գ��գR��FR[��r@F>I=�M�_�:ܧ���S���CC�ww��dX��WZ�Q�8�=C$\�� H9R�S�I�^i��U荌����39��s���`�d�Y]L..�����I���M9lkR�d�������(...`��)�CW��m�����{�߽��Χ�H�N�sǧ�N�0�);�:��^��V�WD�c��������!AduP����zR
Q����a���[y�z��sܫ�A�ժ�0(�I5?)�[��b�eA�X�#��G3-
>�����p&�rJ�o����%ub�$,��Uy9�=���c��׍ǚo�R���]�r�ލ��e��Ӎӭ�0^�/�+�,_7s��e���+X���NzN({2www'��5>e%X~4�d�ڵk���C���G�B�t�������r��囵tu#���x:5##��&2�nF�΃$�n�����R�	��;�ϯ�͢_([4�=�)uGT�D�5<��Y��2���=d�|��2�:�}�Qءgx۵�~�̽��h���ԟ��H�K�����⤻IZB�8y���PEP�c4 Y�N�g���i�j88�E]��9�r�I�]��e�Ϊ撩�Y������婎��ojj��ۘ�lIK�Dw�w���9�&T�,��))0��v�z�j�}͡?W!=\$���57�ܺ<�,��z����	���� �����Xj�F�F��_-����h#���'X�s�,�E֋�-��I?�#  (��Ǔ,�q�9^�֔��/$R��4� ��?6>�*=[�8��&hib�Gxx:��O���M�/�zӭU1��ꇧձ���7d����|�� �`0ã���|ڹl3�֌T����sM���#�&Ï�HK�����T�>���Jܺtqj�آ��G^Jj**��[o�z��y໧�؜r�E���x�!�������\*�XGF����u�A����6QS<�#�w�S}[H�/��YlBn̤�^2$S���B��C)��1I�d*�f-"��ɕ*�nn�<d�S;I�G�W��?��C���z׉�2٨Zl1UϏ�y�˖���HJdu��1�~�rJJ������e0}ю�j�s-�v憾��ٚ�0=���iC5�c��s�bލD��"R^Ϻ{�l�a�S�e��ZFFm�yTO~sdnU0�������0/�����}���v]ASs�y+
�<ON�O��n��0�l�}�Νb�Z9B��x�����H�#�g����S2��5�Ɋ��v?r��*��6�5��7�]m�率�(R
���I��^�"��L����##Y$ڝ�mLVOS0^4Wj-��n�M6*8���k$�7�<5Wz�D*[/�q�n�2�87Ox��S�i2�3�"DFFVs��	���N����d�#y�����kը4�H�f抗�j�f������v��z�M�T�aU8�i����2.:j�*�Q�q�}���r�s������Ʈ�m�����3�v���3�]qBT�,���u�������we�_,3��r��ܦ�ӭ�R�Q�sb\�9"���y���Hj0��jL�3�pv&�\��*aݚ`L�%^�M��Ή:�}p!�cl�K?�K��z���s��݊�á����J����P}��{0���ȸ�UR�ŷ�o���p5���T�?xP������s�[ �	2��u�̦zXdm�e]n����S{� x?�Qov!��2�|QؒD��"����A,
�I�cJvuR?@P^�o�娭0?�(.���������Q�˟�7�
O�QM�A�Ņ0���  rST�:�<̿�8����:��CWW�e��ݟ��+�;�N�ZGRx��E!I���f1�����8��Dq"!����[~�U�$lb'�@�G����d�E�����6R������pȆ�|n=]BWH%�T�3�i������c�+_~�B6z�T�Unn��p����!2B���7m"z<�����s����!������{8��B����qo�06����ʹ_3:������'r�Xt���39��������*���,����o8:�؟8~�833��ww+���1oxsO�03��(�K�����'����E�s�.�aY�DJ���0v���q���R�Xk:���E��
����Z�0���>��uuu!O�x���C�^~����CA�]��@0�c�Ν;�&���{<�<D�@�7g�̰�9b�ޠ��q����!��͂����Ό�����h���w�bcy�N=���4�y0h�|�8a/�&�]a�:g�N�g�Йhkk��r�좙�,������i�����A�a|��a�����5�[g~?�OmvCfLsYqA�;s���G>;q�����]߇g��DB"���%���k+t����(]�t�T���Ј��xUp�m�\�E�g�'6������.��/�X==�Wyyʎ�ӟ{ݿ���d;� )���l-f�>+�����7����&1��l����x䞟g'�$2��0*��߆ey./��zz��%:�EǸپ�������,-���{aK�"M<f?��Q>��+IL����\�_SIM��s��21I3&���	�5�k0�]�}��Μ��l�UU	�g����($QV�V���rc�D���e"� ���C~ʒ��9�����)�&9En㘟��>?U	����8�:Ɇ}��Ri��Rdew��.�ˈU��n��e`����R�0_	����x"ɴ?�|��W/�����D���?��������uH�x3�\�qDD�����d ��$��pH�Kٍ^����ۇK歁1I��ޯ�v],K�}��+W|��� ��4���R����"��=��T�/�c��JKw�,u�tR��x�= lX����:�S���qpp@���o���!������C������B��0>u���OK�`����g����CȻo[{l6646Vf��{H��<�����{xc�	gE�K`u�_z�B�i���� �:!�Q����W`�3�ی���K	�pهG��A�K����yB��dŞǸ�?׊CA8��:��y�����If�ux-==0��X?�Ą�}��c�g��j9���K����(���"��Pd �J�7ݺ�-_:ܧ� ����i��J�����1���QA�)��֛}yuUԼ*�yZ��u����I[D���=d<M`�Qu�c[�w�;85�q�d�{���YH:Y�c)���y�� �m��D�:�aT\��U�vr�%%�ggg�}�l�����L[_�˗��)$EԄn�gI3sUm#�]���,�H�H��,]�Ƣv�d�A���	�b<
5��.����a�v_�kQM���H�ud����,�Ůĥk���B�� cCCN4����CYכ��J�Q���eܨA��K����Z�UZ�|�tqq1�(qGN��c!�p��˾��E産C��* ������C��������<OM�X��rnG�M{��--QMM����

(�!���i����Ec���5z�4J~rʹ�͒:|$�{㓔���N�с#xo\z�!�6�
T��9�5���0��7nެ)�+�N�%o����EJ���XOm����]<��QP.��^9���խe��5ݱ%%r�܊�u�����:�RN��'��2p���+KaBa)�%�\�����p봸�=�B�� �����cW�C�Ҝ�e��l�P��"i�o?�������/I�����,��T�<".�X�p�һp���*U'�Դ�ۉ�B���כ�oF��	%]�H`>~���F��k�ޥK���^�I�̴���Q�%e�uأ�*J],��2�����~u��q�Z�_#��X�Yu�Ȣ@R�}��C�/@�qF�:Ec�k�׈|G=I����G�Xl�y�:2:wZ�Y�*�Cð9�PL�٨g���"��|��B�!�Y1��u2vB����lVgz^�?�'X�9HX,:nϏ�Rvo�tyz9��u:zqF]&w,���|"�uzz:��ӷ;,�3/ف�4
aꋥ��X7���"/��?�`��� �mY��I�F�ʻ�ө�%XHgz1��3C<�z=�������M�/n[#��%�$"n��j�kew^�������X�#��v��8��V��WM�=J:_s���ANV�;��y���>-/.��h�B'�)�� p�t�7գn�UsK����)6LLlv�*��̘M��&;��]��		␨�
�0��aW�.Q�Y�'�6Qc%�L1R�V�ER�6��������CB�d��|с�=C&gg��z�y�������I�A;H�(���r
O�y��	�0l�u�R��:��P+P��_-~�����"ؙ���|�׾mmmZ999Z�f rv��͞�/�a��uV���)@4���.]\@�9����q���]ee7He�3�l��
�uR��������0d�h�����_��}�Ơ~-c�����7n܈����>w�-U/3x��Y��8�h��:.�#~^�ok��ez�L	.��+�7�@��E�ĹI�h+2=���tq�!����+���#��0��]J�?�vHFN�d`ˈ(��T?�4�Ƅ�ֲc�5݈-�d�3�e�"j��J5dv:���$g�"�k���X�p5�,�Z��X�:��!;��͌ҥ9h!x{ZA�C��ސ�ɫ��=hX���%j�	斏Ʈ󉘛���s,َ҉�K㨬�J��F&` �o�s	��Zbe;Y_"d���@�b�Q��0��:Z����An6
2t=O�?JC��I1�Vw+�pJn�l�BMZ���v
�M����$ J7Wo���_���O�>m#�Nʀ��	�M]`M���|��nSDqy����%J5E�2���>��@��Ȣ�=�*�]����_� ��^ֶXq�W$���n��⼁�6���ظE-�Pԉԙ��:`���[YŕBvq����i�<�6:1q�yd��h5�/�Y�<.��Њk6B3n���Y�܌��4 #�:P�hԺ��Mi�L���<�q���[�W��ᦦ��K�e5b;����~�'ʦ
�5�<8���=�AR����P���T��ػ�xzQ�o�֬d��)oɳ1�׸�;�jD��

��أcccr]�0���);˼鸹��� K?E�Lx�9�=��Y�bH��4Bg@�Y}~�����B"��ZO����w�ޤ���j {"k4n]H �Ine�,;	�� B�{ooRm���uxHˍqYwV��`�%3_��гx��FXP?�ۛ�+�%�q����e�Da��z�~t/��L���5�3��>�wtǎLL�[Z7m�LZu�1�k�5,������wd�������)bB���Q�$�~��%����LiN@���^!v@��-��ء�84�;w ��>�F�������Ɣ
:�������/�Ə��r�V2#�H�5H��m������ˋZ��[��x+��g��>e�v$=�8Ib<!�-&&-�:���у^ޖ���G�/Z�63%��R̓�!Z�k��P"{�ñ�4�i�g�S����M5�jt+@�7蜭
9���D�.y���A��ao!�L��|�F.s�D���F�!ȓ�N0VfzL�J:�����B�l`�]w�p�}S�����4�KD�����3ޯ�9F>�A�鐺�ΟgG D������Hۖ��"�qi{����܍�!��jnOv�Yt�?�)w���|"�kvv69le���������q��v ����C ���}�D��0!�v�x"� L�����cb��Y�/�yu�㶈x!>Li�y��%RY�Wx��h�'
�;��Jĥ�
�}���:�Aڣ�`faIҠ�95�2�n�4��ЗH����B��WWø_z����iS4�ĉ�q�r���u�+D��s��c�A����h�KK5<�D�^�=��z�OK�}�UIVbGC�	��r0*3�b�QY�wɲsHX�����TV�Qؕ�Sͣ��U!�]����Ͷ��~?�v���� n����d�P�̑n�g#j����2�d`SI�(��f��o�*�ink�B�r2��܂۶����,&n�M�,��Oǰ���k=���'�gGa蟀�.�vUT��&��X&u��y
<y�%yR��T����VN�}����P�1�1k%�|��46�ST�:V/��ǔA�A$j����2�QZ�&ɁFl��¾f��#�)u��i��K�;�Az6��:�*3�7�<�;�`;3���Y�s���uA(�v	��4�=8�ʾ��>Dn�
j�E)`�|���!Sh8��X����hD���
p�����g6 g�����J�(�k,֑�{�&���e#�HQ���u�� ̻0 �E*1��1��Sh}�wt 5S���q��t��]�J���cSRP��WŸ����	f�:��G�4���_鲐�?j�꓏��L��Gb�uO�\���r�M�)ӄ;D~�	5N��A:�����M��yT��ma�sLj��&�zz���Q��6G� 	4����MN;`"~ZqJ	+<^�r��x�����/���9�pw�qP��{����сO~�AjMMMX�\YSSs���ԗ{����)w*@
Tz��ڰr�R&�K֔�ԑ��fj�DĶ��3J��p��'"��l�q�`�P�|��G�^�H�d�б����ZU{������~&�J��2#���6����S	{'d���?�mi-�#��K���'V�>H23�ۨ����a��l7��DDDh�=����b�Ce1�}��0���^)�G�<fPhݼI�h6rL�Ja��xuW��.��Y"j ��x��2�6J���>)�gQ�V����r�w~�T>צ#����#i�D~���¼���x���w�O�Q�d�Mu{�+���,W�r*H>�� 3��c����
�XY���� �{
X��=�����f`���E� �@�.��$�5�]�TUo����FY��o���Q~�va,��&��<+K5G�rf�vr�{E�� Z���=n-���RSfT��g��!��j�	ʚ~�l
W�a(^ڱ
u١z� ���' �6œgQ���y+`k` ;�F_���񩪪�<��"%kc����Q
�)dط��χ�n�`ع��.��Q�8�8ر�hW���@����
�e_v�
�?�L5�vG��kg��p<b�O�W��5OhSxx�o�F��V�\���<=]Ok�
�k6�S���yFF0%˰Ə��B�^\>dH�=>�j:�q���.�	�̽�>�*�PB��ѫ�L��x��k&�L��O������Φ8�����w�i��<`�8�pSF���/y���Ѩ�J����J:�]<���,���x��×�1n�ŭZ�������A6E<Q2�j��u�O��h��J6�z݋���ݫ(�zO�/�/44�R0�����~=pP�hkadHU�`�Al��Q�*�}  5�+?~\GWm��JFb��BC�Y�.���MX���H9P
����<�XEy7n�hV��Ի��ⅈ���PH����%�S_Q��TJO���u��c�GG���2?(�ߐ�bE��-v�{B/ 2�L��'�]F�`D Ea��2S��pT�Ӕ�����X�3�J�c�~�@�0>E� �P�?<\���������I[J[ZX;��:��DT���C��@@S�%��9�`۲��Rۦ[4V
�	`p�H�VN�<ʘ��{'��c���^�խ���GU_�{::6\��H�L|]4}:������G^�.�8+7��r#�1�݉���ʼ<�D��^^�޻uF�{K�X�	/�L�?�ޏH$�IqE@n�G��!���M��	����&�o�ܼO����u���_�%��q�������$��x�Ow�����W����W�&j�VN@��WX�踞����U�c�8�>0���@�w�ct������7��9�\D��r~o4+$��kAlv�/.D	�E2�hyxx��O-����Yv�T266FZ�1�V@�9�3����&��J��L����IO��5ݔbP����7�����=��8n��-��̓���Pj��l@�Z(��쪁�ch�V������\�h���իW�5Rvya|�8��s�6� �r�Yݒeny�By E��>���V$G�]6�S6]�˽˜ঈp��21}�j�@.�N��Ać����ς���AG�a|�'�ƨ| �>�J~S.)��%��6U��ڿ���OQ�r��Uកg�cD���GI�C8P��P�/Û�/E��s�{�h��c�!v��v�#�N�b�@�no�֜@��9v�9�퓀��� )G5�3�ފ �Da��_���9swf�t�R>�'�)�R*�6���sb����

����&@Q ��8���Vn�X��(K��]@5���mG�g�q���b�{{�o��d��.���uG�ЅW��U��ܞ�,�Lj�B���Z�ῐ�?G'�ھ�\������K�X�k�`���8\%Z;�C�䂚�>�4ee����>�9�X0&$$��=cg����߁�{������î�9��2�{���k� �)W��mu���z)))�0�e0�@�����.��b�e��H��b�d*'Sѣ�O�Ao���	���򳪨���AU�njlA�˛�e\B��_R$0G�k�˱I2�ߡ��+66���VA`y�⎺��.�ꜳ��4�ѥ$t��.n�ߣ�c���:�N�����A���E+� ��S�n�r�b4����K~�3=���/�aFU�ъ��r��-���Ы���n�1�}�|�5���"��Kl>�a#�YhnnyIm |����*t�1E�'�r�x��ȆXH�����B��:thT�sB�w���K�_����
��BB��@���kx�.��R��U�:�mܺ8Љ5d˹���FFF��Þ?��7�.F�����(�FA��ϔS�v��E���U���@G0ԯ� �> ы
��7���6̼��t�ċ��g[��:��k��:Ŷ�J�Y��}���c���'��A��{��7����X	���`0��l�T�%F�P�̼�+1��r��,�T	��-,,�����A�:�42 ��뼎?��9����D��FQnq>�f%���*U�"��|��^��Hq��Rί��ji1�:������L�H�Ofz��<QX��Zzzz�ʅ�y����M���?%��m� ���x46fO�H�\�~ݰ��W/ �(�4Y�4�F?Iыq_����1R���葘E8";c�04�>�+��b��s6ғmvvivew��b�0�ʓw��#���~y	�{86�����u<	>��m����7���}jh�7�l�A�e�V)�#�}�Qt�k�&v�=8�SD04�vw5�.�ܖ�;BJjJo���)'�`����!%�ݽ���=�-��9(���!yd��X�mص#�t&����A�������#�fdϛ�麻���3�S�x�Q���/�H�dmS��wWh+ڦW��]�G6EGI�帖���	啃dr���<2Y����x�	:GV> èV�N��O�H�.3 <ѹ���Tp�'ORΙ72��+sEEE3z��~9�{<��|�$�*UYY��-�t��v�Ζ;��={v�g+qT�L*{�P_��y�a����.�O��	����vS.T��]:�A,�F�NR��qv����xI����r��1���(�u��;�v,�Dw.�����R�b����u����F�G�tK�T�~ѣծ�(��EҖ�����T�/}@Q$��m��eSZ���[� ��3H��H"�4+��.Q��7��
���@����PzKQ���1~aa	ۻ�#���ZN�m5�!��"�G;�
��tZ��_�Գ���w'̍� X/�.N�#�~/a`�N����εs~,�pٍ����j��Cg�讽����\�h�M�A��x'�1\@���	�᪞����Ћ˒���9���&Ƃ~BGP+WFD� :����o� h!R�{�-�#@� F�Q��;�y�P�Z�����D�|�AO�O׊SB��(����h<@}��8nE`li�s~�&3`�_//N+�R��m@���*��U�X�6b%�t:�%5袞��(� �#����r�Z����Zq�P��?�\2}��f9���.��_	���� ըe+����aJ� �|萐xc������G`�T`���0
��T�^�F��������o/�ɀv.G�G�d��?{I�V����ۇ+~��5$�P�<�H^����;v��>`f=��y_y��=B�� `������/z�:���9�Ά]��Մ��Jщ2���gm�	L����pr$����+��%(F�,6����Fm��@�mQ��gՌ�5�/���rFyN$���#@����]j&sg(L��%�&����Ǧ���u�?QeeT��1X���X:�Z�o�������Wj�i�{�Y�~���F[�AZ/����A�:y���C�����Qy�H�cS��y�."��}}}*����$D�������s#<��EZ�����sM�.);��:�D���υ���7I/we��w����G�~�U�c6��~<��z����6��ƛ��C�~Dg���4v�Q[{_�?�o|4�{�y��硭���S=�Mt������M8�Ǎ��$�bZ����Bx]�#��~�ć����D�v;;,�@E�;�x���{"�o3���'c|��i6��&�z��<ʽ���1D|���v�m~}���x��4mL+/�-��k�>f)B�|�� p�E�W�kʼ.?K����$�U-w�����b{'DnNE��Ћ:,�Ѧ��e�Ś҅ {�t�3 *yDA�Mt,/v����Р�ݤ�A�:��������4��*�/��K��%�i�2��өO��a�F�|9���J�Erl:�ҍ��`���:v��A�K?}�">�%����*��!�O1Nk�#�z��{��$3���[�][ڑ�O�A�loLs8�v��L�D0�4$�h@�4��9jO> �]m�����R �#-��E�Ν;MR���ӂ��0�@1����f=�]y4#�X	t�ϳ����������N)(����wov��=qx9�/��z��z��Lt���Pey:�+A1`����s�Nx<Y C�;��[`f�1�z�oo�3���[�n.]�Z�_2O���vb�K
�c���=77��z��_�}�?�؎���������7)������dքH�kld�ϵ�l��!m���Dz
lW7(8�|�1��dV
��޾ͪ{�1*B�288X�UN��X�Ɣ��'�;��Y��_i�ndccs��l1ǽ�o��.O�}������b��6��dv5[f'��2�ij6�2N��=Ϟg_�s���\�	~=�����Uv�ų=QX�@8�䙇r���ɲ�ȹ�?����SH���`fjqqvm�ŋ�5��;�|���v-??�e����� s�˗�X&i"[�]%L�o�Wx�}�I��f�~�z¥/i��p�I���/*xΔs�1�Ӓ�h�lIe4׿�z�-o*�������#���XmC�O�.RU5N���cץ4�Ь��V�Y0�Ž���n�x|zZ��A������w��}���1K���$�o��6E�>��Yv�R=}ݑ&g���q�o���F���4"�Y���N���;�g�����t�u�>ncF�ǲ���Mh_�d���Zi�N�cRJ�6����r~����hwUa�89R3KR�^��5biɣ�9;G��] �@d�B���Ǘ𷈤+<��		��z��uz���Tp@Ȳ��^$�_p�M�q�����+7��k ��q�^DH���"�W�KZ\\<���U}qq��?�h"�b`qM��`zZ��E�_��20�@�ƺ-�/�l&&n,�T�����j�AG~u��器�y*�s���z;]̰�w���XŹ$Ϲ�ꏏ�Ů3�R_K�Ù����O&���rȮF�ib��bbڈd���ߒ�T��0� A����0�q�ܚS4� 4ū�M�:Q~l֭I
� �4ИFdgA��$rt�G�BGC<u.�ᇆ��v¸p����]�9�H�8����X�5��	���8d��[��~�M�W ۀ�����&6�RFaa��/��7��/H��T��񦦦^M�8�M�~Ih�J�d����g�ݡ�Hh���a��{id��~�̅ό=f/��c��u�v��,�2���O㴍αL�%n�E�a�m���H�� ��{�f'����L1��I�s.���|� ��F��}dL���kW�f�ad���Y��q���a�4��=F7�?�d�dD����)A7;vip��1�Gn�DwTB����x
���j��2զ!�tI΍�,��&2�i�,�D���v�Y�ﱕ� �O�m��`[��ۅ�Y��YJ�=�\Br�*0�<p�|������iڶw	��z �%pΗq�mhh�K�K��Y�	@Jj zL�]�t	�a���		��tth1s���!'MLb	�,g�TPp�(7���Q
.B�LG3�u�oJ;g[@��DY��=ʯ��o2��	]n���S}=�j�;��e+%i��Ra�w��v���F����J��C��!���l�!j���:�O,�2�������۷��-����I��)�v�~�)��1��w�d2�����V/���8$Z�̛�2��x��֕I>:|��ev6��M��D���9::�&�c��I[X�8�Q���){��T�cWY�ʮ^b����� �ޕ����I1M����o�U%���y{��� �y�<~�Kέ[~���ӷ����@2�yp����7LT.����_D*�D��g.���~�g����1S<���)[���0}�����e�m�[���P��8~�̀.I����#22VT���	���132�6Gv,M}����*�㘽~�}VZ:]�+CEL0�H�qƽ��T�S�y�i!��|Ȥ��*�v�â~�d�ê�<{�ۣ�v����{�fY�@�eѭ�[d�u�s�1�,�\���ڎR�[����|��K~��xmmm����ׯ�2*�	����L���{	�a��5i�1����i���*��m��~�E��o���?iz�m�}(Z�]���CZ*#]e/���I��G2� v�DS^I�2�{�n��ӧ�B@�R�����9u
�=�Y�1ʦ�^��IH��D������Z����x�@�]iLѥZ�ʅ(	��o�w����4���^�{�QUS�>~�G�e0�V��5U,���6�i@��[�ݧvĢ�s��UP@���.h���տ��p+��!��	w�ڵ��a�%�ג@�#�d�t����2��2}?~���ƀ���`~Y�i-�)�7@�&��Wo�VE�[��J��6t@�����yрf��e~7x��5<M<��=h�{��ly+���t��� =��mbB��6��(��~&�g��
�.�=>��m��}l�s�Ƥem׿��"��pJ>ML�dp������Qq�%�����@��l�/�۰xy�v*��ZXh@!�w:;�����8����1����f�{IK�hJ��˄����z���'A�׼���OHH~�ܪ�ȷ��e�G^�d0n�Fd��.��7��l��عs I~1���ð
��{Eh�@F UW�Ux��4NG��A(��[M�X�Ƀ̄����Y^��-�J%A�U�jy��t���x�c��`��,��bbaa Ȥ-����|�P>Y�r�wö-ws �r1��3��z3��у&%�����������k8)H��Ѯ�q]�K�0�ͳ�9@�x����`��V�@����QU]@P0��+ `!���}���?��4Uo?P5���b��Y`�ɘЯ��H⹊�\�^�*��x.!!a�J���&���
�A����EkUqpȖ[�1���/z�1�"�b��?����a� �����{6��*�����}��s�U�h(��0F�p�V�\u{u��o���ÿ]�_�����?M����2,M�ѵ_�_Q��jaٜ����(0�9>�q~��zLI��_1L`DoJV�G*�T5��%��F(�'Ҝ�&���Ǯ闸�g�&��'�I"���_��6t�c��q��*?Y��+�Y{ěVYhY��q�s�˰��ΝsY�퍸��6�[o%J�HJ>oLՃt�
�G$�l��3��/$B��%���dΓ315�ĸ�7<�t��Oi1X��Y>$���V4���2�)�UG��I��ЍQO^�� AW~��.+�e��a�n@���/.��B�`�QWW����؀fF�Rwlp�x���j���d�
Y���,�b���l�C��끙'�g�<���3O������qtI��6+���~�p�Sa���{�8l��r���u2gv�����������-Tɚ�*�7ک8� �}�Qf<vd=H�4���T�#7�#� �+]�a��v�ݻwG��d؛���$ &VP"���4��*M�R�����87	_��X'Z�}�į�l���1�O��t,@��x��n�s�Nѹ@��z�h���>��$R��jH�;}�=�Nd<dy&dŉN�l�]�	�hT�.:G��a�Kc���a�g���Z��M��g�StS��Q=�w��irLW@@��M�������D3Z!;�J�Yy�U+AV���I��s������g��	��m*�A�]�e�s���X������Ů�����֛�S�>���;�ž�J�TDYCZP�d	�-�ز�Ѧ��&Y����-�#�R�PG�Ph!��?���������u�y���y��k��~fZ���<�3�kr���T��l;��o��ߏ��Ղ�������0�枚˙F�O_�U� x�V��RV�	.6/9�	>�G�IJZ�@��xɋ��o�u��3��sѬf�?a�����^!�����	׃���ij���U�x�C���9oE?y��*�0l�t��/7���Q`ᓮ{>��d}Xe^DI�a3$���dZ~�:FY�#�W�/���나P�[����4��#_r��N��S[���%-��[��%�o=�{��?m��9���ϐ$Y�G���{���;�������7�+N慞)�����)����c���p����D���GC+׮�{�ҵk0��6E+�b.b��Cs5/~$��[,d�C/v������k��}W�k����ۖ�R�:��s�������*z�}�^B�IFY(�F]?�n�rt����O.���0[�ߦJ���mlh�˺<==<W���(�꡸@�U�菋7_b~"��6�RG������$\��+��~Z�IT���I�T|����<>O$w23�s�, H0l�Ѩn�A�Ӥ�sqr�}41�:X�+6��G̷��޵.�"u���6M�z�bbu�E�n���ih,���>!���ϗ\v�065�-������}�����5;"�Xk�jr�__LMҜ.R�r�|�s#�H�<s����n[�+8�� �yp%�p��Ƒ+�J��K�#�:r��������lB�˺�;s?8����	��<��҃׭(��~,ή05���D�.�s�� 8�X�_��Xtf+>���ߴ��G�
����_��;�z��Y��	�(�G��T���F-����)��]�&:r�����p��j����@�����2w�-#��ѭ���.���5###f�����k>�_!W��K-U;��3`�~��#�_��|Ω�':8,C�

6@���E��R>�[��f�9V��Q?��adj��7L�[[gc�r��f�_�2���O��5����P�����毚���/�6��u���=���Ϫ���FjEDD�����0���NP[��� ���r�y�,�����.����b4\�|�l�3���;fo������4��l�k�wo�<GG�)��l$<���?��9�
y��@IR�������߇r'�����gՍ�����\Z�J�Pk���0��nnYR	��$6AN���~�Q�
����u;���]01Ȕ�n��D�7�WR��&=R���m����|�Eꍐ��DB
�0A1���w%�
�*{���H'B<�=<��㋄��Y� �w�}�$����;�\
Cd�Y�[X�||.4�I��d;��m�����r��Z�	)�!�eʆ �x�G��Ā�Ʋ�FT?� I��ם���1�շdZd�<8���م��ѐ���	�˚;�y�����7A��f'������/p����>����ꁘ�����J���LW8/��EQ� ���o߾v���D��4Z(���V�`�R"I�~��_�1�����Ɯ}率K��v��+�ظq��o�}؆UH�M�ɑ�\���Sʁ���:�N��C��g�8�[b�ns�˚4�`�˗{ �H�ϒ� 'w�8�|sG�]>>�$%�֯$�g���i@�?�c���Q�Q�D�qX\�����m���@3�ED�	'l�ܖiII���� 'e#G��ڙ�����GMì�~�{]�,���+���L������\}�w;�����x8N�%�dU��]���Z��3<�			Y҉A��,c���J�>;�{�)|��A«�p��R���o�[�'n�raQ�8'��K����J���V�wy�'�َ�_�*4ݻ��fZ[W�w��(�~�r�����j�A8 �8��V�	~l/<�ui���f�����/����˖�kη��x���gq��#���TY<��b�������\ s`Z����Q��`do��9�/�A�Wo]i��S��*t���*�.����gϟ�|mN �8�����1��������c��LDm���U�.:�D+�����uu��6O�)a�#����a�X��� Rx"T�
y��	ϴ�XS���6���Rk�s�yc9hm=:*i�
!�@xq�������|;����g|�㟜����#7�����Aj!��D��l���9���{���4��:��,8�1�	���zg�;Qc�?67nm�ȫ,��_��U��c�`z�azix�+/�	�t��! Bۥ��J�*�~�T0n��u�~-�ɐ����J�b�iچ@�m�sihmy�|6o���u���E���ʩ%��+�n�1[J|�
�u��*\v���_fuD�8�^��K�46�cW��:�2w�#�����;@k���"��>���;w�Z��ܧ%�B2>��7��M�W�޹��wA�elf�}���\�!�u���#vg7� >ڛ�L˵�$'!ʹU�b�*�N��� ��e�#o]�����+�:�<��'�<��8�v�|�~�j
z�%��� }��/���]����U�Dc}���oQ3���>������.��z���U]g��Y|��E[�e*H��>�Ƈ�ԑ�]�l�Q�>8	:s�|�O��I����~�q�����n򠾎�a�+XT~��'kAjj�*S�л�[��7�u.��J�һ0Ѯ0���<2�⣼�$ �h�����4�Ʋ��<R���1`㕕�w��%OX���������?K������ �/���k��z}ĭ�l��qV���;�*�Sς�j��t"Z�ќӾ�m��� �������#���J.8�������\��odt9��c˖-w��[�����!77ܠ�c&�UC^Y���葿��^齺�DR �~��-����6���L�V�A}�ͭ��*�>|�xhr�ם�,rwVx8�IQGWy������]�bϧ��q*F����QL������CA�v*Y�9�;w�v~~�jy;XS�������	��1V!�;�F����V��^\*��@Bn,��o�"�uiH��\V6��ikk�U����1ɹ�=�P�U���ǻƳ�4f,�	(���3[ݓ:�s��i��	| Jc��ywn߮V�[�:��K��O��|�X�h�Ft?Y���Ĥ4N���y�֌�#�0�S��?
0quu}~��V���Դ�H�W��W�%j"���I���o���|>�tr$;���f;�4���B�DUU�+[�$nܿ�8�H�:��pb<��H	�qrUD2�����O/�[�f)mؐ���*A�;7on��/�����9��L�������M뙳�{+d}����ǊO���+��L�򙚘�R� d������/G��a�7����(������6_Ȇ%��ԜZ2>%��r��A�����2Ѫ<^����l��n<�<���������{V�6�|���Z��Q�%������j���e%m?�;'g�}]�}�ߚ��ys)(%=7��!8���s�'h�N������l�`6�:�q/�էDd?��?Tv���ݻ�G� �W���fw�3�t2�����d}���Kw��	�?̴���?�����k���oK|�!�^�v--.Nt@�VQ�e�Ye�%"����L.,4el��d�fC.���Чh�����L�nMN��Ȫy���߿L�ulP�o�����K����3��O^M��O}�o�2��K����̋�	�&D���kK�o�4���eN��
[p-���M���A�� `���ANsi�r�<l��4ѽ��*�{����k�e�'����ۮ��ד�w�����|}Uל\\�$�qpH��'����/�w�����hbgle������'q� j�AII�w/j�� ���e`�u���6����SQQq'=R�b����7SQ�����	�5��f��~�u�4p]�9)��ش헥��ʖ��~����YS��6�7�����ϱ��2��w�j���in�HJ������`H�����$<��(���|w�K�'��_`���kͥ�0C/�x����C-�d���b���q`sCÍK��ܼ��ug����������g�i �1�!���H�Qx<���9�!c�;������`]"%׳��/^��d�	����[=����/5��B�����o����;�����2g�rI����><�����g�r�����e�VJ-�o����@��Q��c7|8(U�E�>��K��8�X[gǫ������塀�����f��m�%�ȃ��Pu5*��o�}�L`,��o=LJZ��ڊF�|�����I�5�#�!We�RZ?�>M�tUwk��Ϡ-eH�1����+R� ȃ7�⮂z��h�"A_�pA{��pE�ɹP5Øne��[r�j�����'�օ��)g�E��p���[���K6�[�]Zj0h+��u�2D���K��\��耬R�?��N.A�\ED����bbc�8�L��Ib�ǿbժZU�54�?���=�,��$�q�W��	r@�m�)ɋQQ�ǎ1ÓkTY�;�&�����}��SU֢e����0��<�4�z�W��ADt��O�̿.���,����/g>u�.�q��dWГa��OODh+�=1�"�_2���ᑃW�q�瀢� ��[���`�#4b�!i��xzz�v==�ւE�?� ϓ4�9wm���f\�;%�&O1��E�D�܌��GYoW�9 +Y��Ջ� D�Ǝ��*�����ھ8u�FU�B��̭���Ϟ=362JvnJ5s,��$���de�G��R� /Z���m�D^m����-s�	<]�k$����5ı����i��F.M߰u�E�3fy驩�)))xBə�d��9h�!��������̢��b�u,�d*b����f�҅����Up��tnTlr� ,�ML�b���ۼT��#�<n
�x~]�e�N�5k���Ӌ ��7R��b��V�~�������"b�5�IL_g'']���vo�~u��z2�H$������TTT<�L����m�S2������7y��<6+D�]��@�3ٶ�$�q7O�)��<��u��q�j�+�s�?ʆ�Ĩ����w"����EڒP�P��ލ��X|o���9E��L�H��@��,�K|���K�w��?m!߱..B�R �Eݭׯ_��z�~�
�r��I�xR������p�ӈ<E_����08�k<u��K���F��r���t9IP�=Eu���7X 
�Cʻ�?�̑�������y�Gw�cy�g������[UK'N����Ͷ	�(`Ïϟ��i1-���ҷ(t313�ο��6�Fs�q�v�2�8L�V9�+Ʌ����_�ƁO=y�y��{ZW�^%ώ���9�	a�᲻{1y zVƖ�;�h���׫W�RS��V�r8��ڮ~����������ny�֙IK�X>��6����?";v�(�4� ��d)%ʭ�8X!��̥�B��?oߚc%K0-,�R�d�
��ۜh�]^�5`��x6��$��]w��E���RJ᧊t}�y��R���u)�ғφ���������D��b�Tb}h�C���`�-���xYڠ@��Mg�ˑTކw�&�3���vH���k�e �E��;|�i@��׀)"��$��ϫ���\�� �m��'d�xpZ!rsVi����]�G�W�̲e�/�Ф�����׭���a��q�	d�O�C2K�B�°BC�<w�&a34Vœ��"&�0�Z���\,� �=�g_��f>�,�p�Y�PɮY��n�FFgH*���X�\��o���E���G�JnV6���d��ITrK~6GFFa�}�r�����!���\Z9����,,,o�d���FC`VW�\!O�u�Z"�?�\<�$%�;������H;��l"������?u�aA��b�/^p�G�A�� M7�ڌƂ40�/�W�Us
�W���<�=u{���OXy&�3eٵ5���͂(���4Enɴi�2�	��Z�����==N�t���g��Z�ǅi�I���rk F
���;�
%�>-�]Y����`�J~a�E/AY��Qܘ'g��Bۜ��X�����5�,<-Ԥ��A�T����HE�����5Y딕oi+̀���� ��I5]���+B�iw��'�1�=�.Ϻ&���hXg���g�n���y,��7�I������2�U BCZ�����nU�#�R�mʘ�MA�kq��Q>�[�K��a�S!.��򗭯mij*�b��sf�ׯoWVj��� �|������F��qk�	PGk�EN�����\�
�@s HO��L���hl������M�]k��������P,�(e�2>��C�28]�@���b��2��7�<0���rN�<���Y���>>>�(��
�!G��C<�Seպ408���g���e$��gWF�~[��P��y��ё�+��Ő��{���(=9�B�/}�a�����Ԕ!���D؀�z�,�nޢ�����o�ۏ[y���@��٦t6�����
���Bƍ8�бS�[2\_��[_�!: I��c˳n��'Z�� �1��QrO ��6,��o[��,��]��ѣ6"�����W@`�4Uǣᐴ7��W���pOv?>��Ԋ���KT�,F��E1�j(x�U<Z�Қ�|�K��v]L�z���O1�*o�8}����]o�n�0V"�'��B��W$�x� ���
[DeC��k`K+�s6F���~h�;���0bH��CLv�l�ڟA~�@n���C���zc�N�B���ooAp����ת�� �C��J\�0;���W�1�n=�=��b/<� ,fd�|���}-f�h�,���QB*oE�������lr�^p��9��ɉ��!!�DY�Ǐtď�b�t+��j�X�=� < o��X\y3�������*Տ̧�s�6 	*d��m���ԃÎ�ơ��^��Z��E���ڀ�{���OD�V>��}�ˀW>�����9ŏ���;��-����?0�pݬ=�������ON���̿}�Ύ�ܝZXh21`]|�Ӧ��w��'�����zEE�c,Ny�`�ʌ�D�km>����͛7�F�������<�ܲ A�m���[�GL��:�!'\Pa��x��$9rY��Ǐ�̥�R�]�����H���x~8�8�����	&�&��ǿ�9m�nĕk�/+�q*^W���X���?�f�Q���#,$�G[����.����ߗ���x��� �l�:M�<���6$M=!"*�
|�?G2,�.L��	~�W\��#��Sz�L~]#Q12:z1&D�f�+c����m����ݖ��P�N����e��A�x��9r�ѣGQ����7�����!��� ��'!w����|�E�����),�OXke�eKy��z&�ޯ����)a����9��^c���>^j�03�~�����Y�Z�u�l�w.ã�<�ٌؙ>��X�lYuA\�'�r�.#��$�5���������̡Y\�����ލ�g ���� /�2utrbN���2��,�
��y��
�qtt�Cv�����'zS����p�O�h=]a�!��o]'����:_C�4�P�R�v@&݀VM���۠ڐ]ɛ���ޝC���e,�N��N.9��1>����x�(��9Q.�k�B?�m窔�#�dN�W����Ct̗޺m�ggƸ�I҃�W��cR]����Y����|�6�c*��M.8._W������%KT�75>	
�?�iR��l�uy��j_㇂��
Gww���V��_�Sg�'��&����0Ǆ���fkx��y�t�O�V���{��c��_�{�Gz'>�hzz��l��,m4}�@�S:�Is���~�]q�?/�A�E�)���J��}�O�##��Iˈ��ѹ�lm�b�~�C��{_��J|���9c+Z��%�i��2�{ڃ������X����`B��TI�DV�5�u��IB�E�����x�~~�J(2���6Ѥ9a�]ݱ47]��)\��Pk #` [�[��m��X�sj�g7���&����/�����/�Z+Y|���<e������S�X�Z���H�W�<��D,}�?]��BԘM���!�ZQ���|+�b���j?�d������H�Bk9-?'�9�������A�)�i;�V9�4�g��QOu��Dk`���?�S���a��^�|)(.~; EٛNkN�`�_���A�Xק��Goc�CL����u���sm�������Z\�e�ݿ����`���X�ï;;�s�lx
N�yf���_e���Oה֯���-�
d�������� �0L"2����ã�Ѷ�X�뻡`%l�����p���*,���ӏS>@�ߢ@� eQw���i%��,�2�a���Ԛ�~���q�w�K�v``�8�A�W��SwRۑ���<��to�av}J؛��2���S�/�!�v#􌤙,�o����1�TG�J���[s��4r$�N���_�C�b�)fMg���^)P��H�'��3gμ�Kh�8ƨ2B�a"�\��q�RҤEq9 N��Thm��e!�|����Z��^S/�lw�f�9ƃ"*�`��ttt�p�\bx!۠�*��g���?c�|MP/|��G$���g#ӵ
�w�Oj�k��⍱����L��ze<���\Ƭ�E�k�A�arH���;�0�i����Jh�qQU3�=˨\8�i�$}���Y&��^"����$o�����=�j%�qH1�`o5��|�k��^�>uU�̯*e��R��1�VvEU뤞cL"e�{%�&�~�)�C8>{�g`&l ���5I�i�Dԙ��?2�'{d�w�~�p��b�rFk�l�	Z��xç������a<U(n*�o$M�+>��1�Y��E��
�������+��d2��`sxC�Ŗ�xC䎔K�Ҹ����5�.�C�N�! ̍Т�B�c�A�l$,�,��$�kAK,�Ԉ:_h�y�I	�ʒ]s�@�rӜ����+�LYմ�v�D�W7�� -U^���K���"8���tV��"N���rD����_�`w0݄�V:�o������2��;	j�`+�ǵ�+8����c�/YZ���rB��Z�K�~���lD\kK?6jR��k����+=f-�6���JX
4p�?~�������6t}7�\&��� ��y��t���U�u�����? ���*���c�W��v�^R����*��=���c�ب{��;����b.ChNl-��ݔ�j��f�y&�YTJ<�
v��݁�{��3*� ��'s/���$_Vq����O�J(��X�OIS�8�����L�̌ցt��fc�IA�"m:^6�(�ƎrbA,̚�č�uww���`�噱;v<����bߵ�)uԌu�ηč��;�_he8�"δ|f�ɋ�f����R����O,��b��F�ϬQ���O�$ު�`����w+�SZi�&("�t�g����GP6j���q�ꆏ����U�!0J��Э�:� F2�Ak@XPPwz˷��al1�3�d����{U����*�|�yl�ڋ'�}��,��̽�V�iӇ���<����P�+!� *>!!aŵZ��죔C֫��"�g���se}�,y`2ҵ�����♈繬��ò߉|�z�I[�*e0��!�ρl�����#�x��9���Ǝ��Z���%�i0i| ڕ���gdx9I��Z	E~��Z43�n%k��M��+ ^��9i�)��0���/��7Nb��0gAmijk�~�05xh�J����ʊ u�O �H�1�	=`�~��4W�:� ��Ev%{�7��f�q]k*�m@` �<�:ᒃ<d�Y�$Bn������y��'�����-^�v��j����iXrk��e��=��
�k_kA�� �mDg���Ֆ���T���Q���szPU�P̫nn7�����j�� $:se�LO,|۫�p�4Y9J���e�5�ˮ�=�t��qF�LWc=Ǿ�Rt��k�[::��	�!���	�2�s�f���zHVn�Q ؙ�r��(�<�c��=���,��		��A�,Y��bG��=?<��b=g�;�"��I+��vދg&2Ņ��LZ�>��:h���R�T�5��ʎ����9�Zq�:{oFL���Q��kK����G|[U��3����'�V�E��^o��]�yA����%��ep���~���5�"w&�xn��BEM�*++��*���++�t���>���V
[�����hG}N� �Vj�����s��s��/�z��j�ÇeQ~z3�MßBBBH�Q�aXB�(D�|���O��fDb����[?O��f�w�t)0�mϋ�V�ӊ�kxѓ���H�jg���2_H�!,"��c�e�Z[ooE�v^_�g�Y�T3�2}�:|7v��3��@^�����=�v��L~Fp�nan;��CCC�߸���p�m�ņ�Xu�׊	5y�dZ\�Q�ˀz�>4r'Y� w�0���3)���G�	�/�w���[����@��C�5,��Y����&@��z *˴�/~��y׌�v�2�:�`%4=
!�n����*B1�g�e�/Tg��B������Z�`/mpk����[�2��G�P��B �~�h~x���S$W���p��niQrĕ�����x��`;v�	�����C�3 �;���.�"���'ѠNV1�&l˱����{��9�^gpd��n�
x�	v�gcg���};��w��ࣤr�\��<U [��qq��a,�����a5u�ŦB���8����f�6�L��s���
��7��2��71�N;ԝ�?bk�Hql���X����ʈ�6��z��1'D���;�V[ j�A���ͳ�|{��`t,����l��c��y�dD!�Hp�������f�n�� �/ 
����b�NZ�n3�l�Ś���euQ�e�h��(a�� E�Xy��5̀}���P���B��c{�����'�	`�T�8$�?�c#�S\a`��5vAA�@��Ǿm��a&��1�م�J0C��K�9ۻX�c��H�ӟF���&B1
���n�ʳ��c���J'��B����GRٺhZ��:~��)�
�]�v�3R�ՙ`u�m3V�x����H9,�k��5Z�FZ,�a5���dBA6g�.��
�#Y�[�}^�q��:���r��)'!��������������h,܊�Ϝp����#Ǿ6
����� �+��mutt�F��8���
��3N�f��Ԩe�>���J6Lr�s_���M�'�Q�2W�73��P.NNl�����V���?'��m�"T^^����P�XvycE�ɪ����Su�Ũt�D�`�&^��+�Z�m�\FPo�&qU��xFб�_=ܟ6�`T����us�l��6Fm����𺀾xx÷]ha��?ݓ�̫�n���׶��`����Y�8�aI����ྰ���4[q��W���mٙ!O	[��N�FZ�v�e81�����Y��1ܻ�^��r�����S��p)l�3+���dyE�+p����w%���U��e

��p��S��l�f>l��	+�Y��R�"��:!�F�)�k���:)Ǳ���������m�j�m�J��l&"�>M��}�7


�9$H�:�P�0Ya�S�	mq�E�v&� ���h­�z�X�j�n$�H�	 v2V�D"Jjj{��5�gī���Q[��K��	�w�bo�>Lb�����`���-+�$��ͪ��zS�-�?��FivNN+๊�؁�FӚ[�v�;+ 0<8�B��=aIm��_�JN;����:��h��Q�'#D��ɐ��&&O��hT����tEEE^P$JX 9\dL;M�Kd���K���1pF+r[�#���-w�x��M<S@��j���Ә!}U@7�:8)��4�b7�(����h-� >�	����qk�oΰ;xP҇Mq`d�K�]�^y��x�����HL8�Cv]	Ђ�i�s+�A�A��@�1�n�2�<�(�ܵ�e)j�ۇZ#G�r�D�r��-"���s��It��֩�
3X�g�uWyn$	��-t�f���>�$�\8c��~�������]Re>��~+))	{�!��߀Φ#*cl��=}���6WVc�� ��zʎ��DO
;�Y�oӶ����^�0�3����\�|�5�_	5P8������#�z.��g�C*~��Q�?�O���z�G6>�j�bK����B;ʽ��j@��A���:���wz�Z�0x�౮CT�vtt�ąr�؛\�) o�'l��
���[ɗ�}��ϨU�iǣ@�{	`�
Vl�	��AV-�qr3vnę3yY��O�3�-H����w�X vU=��j�	Uە�6	��D�$N�H�՗��9�a�i\� H. �,  �)��F3�s���&̟a��֬��7ia׆-��w� ���ᪧ-v�255��&���1:�G�V�����ؘn0�������(�t�]`H���y�&Ҭ�E_�~�Ƃ��틲��oJ� �[R�b�GY�����ts�����oǦ�e"s�>+�9Q�f����23�!�J;BJL	�i��s�:��O�GV3��2��`$�r���*�p+�T�еȥB�KԚ��d����x�!�`j������!�1�
�>0,/�1��896ޫ)~�X�ts��������lق��Ţ�$S�2��=fv�����h�M� ��p��1�M=�4Y	�WX����㕭h����#��:2:px�k����o< �E�&ȭ��dLz50��72*D�W�+�H'z7�O��E!�׮i),�b���|ћ��%Nd�(�X�N;	~�_����뜕����1p���se������ p��h�އ�v����|�+\zޖ�oW<�^-��D���M�H[?��f�j0�zS�~��j�� rlu)��%,B��='����ַA���3�B�Ug����?��9����g����I4'�+	�ɣG�<����y����K�������1֘xm�w��_p��ޓ�w��h� � M�¾�I k��l�VN��� ;����	���y�=���f��MMN�+H(�ps��ϟ�c��u���h�1�1$�"���Ò�3S�C��<�b���������ua�	�cJ���t���ߐ��ERHHֻ����̹}�������3G�?oq�qf��@�1H����q}�z·�)�f�8�^i/��`:6��U���-5�6��&�/���X8ۓ6���X�ct�f1�-ja��%%�w�=ִH*����uv6B4���L:d`F=}cA��	~���$����u;��,Ì��pw◥����5�m�g���`R��NΜ�����dQ��(al�c�]��y��ͫ��g8
���� mX3~=}�t��A/y9�HU���»Ӎ�b�Ep' rs-,�����Ƈ�Z[����%��vN��~����R�2������T⹨�	�����ۃ����z�!G٨��:|��,���0e�?�5E��΀�0��\�����y��11���1�g6bbD��-����d���0B�9h�o=�D�fv�Z���X�{��(��\kjs�����䛃PY��.����w�4���=���Z������([:�}<6��>������[�Ӵ��E���b�J��oP��$��Bü�R&�+^�޽{�>}��~��݃f���۞Ţ��1_��El�η3�%�}��+��"���tɕB"�{��tV�<g�s�;� �N��7��k�}�.읁�M1�ZI�<�������V�'��1�71�#� ay�Ϫ�132��`s���^/[Z JP� �D��s��@L��K��},�o���g39���j'���q!!�3�A`pաء��u�ò�,I�!�T^\���I�Ý!���o�r��X}�֍3Ww���(�D7s"��F�����[���#���ۀ��8�h�J�G��UL�HtF:�4"D�	�� ,�e�����\YlɊ��go�6���q�ĈpZ�s0TAHÆέr�56�	Wc�p�3�Ȼ<
�kc��ao)�O>l��,��g��e[��A�l����ӊg�}	�]P�<�Ӳ� �:��e���$�6�sr����IWά�9V��<0����z���åd�}`��އ'�f⪦-�����F��J�Uf-f;;�AV��|�u�aXƙ{�S�Y����z��f��"�X�Ǽ�`V�� ��:��^��b�!���b�i6�����cSv�#B�p�<8�mH��i�賰��5׌�-Lk�J���^����Q�9����ʊ�l�Ӂv�}�V�y���$'� �ʏ��(.l�bx&Y�����Ǻ°�i�5G ���ʿ��B����`_Zƽ��2��_�V��T��hF��ꂚG��t��ޕĮd`�ب�\:�>�xrrrү/��M�t��M��z�?o�!�f]U�Ob���0��߅A�������bj�w_�r���Ǚ�̫�@� �֊��K�ut�O
X�&�m�' q�&E��ܩ��P���^s�!+{�p�ģ8X�̜���6�3����2���@'d�>�#�9՚J���{�d[�]����gk8'�1@H�!<�Z,�#�Q �i�q�/z�����ζ�h��|�x��V)\w�a�2�y�=���X��b��ꆆ�$4ҍaTJ `s�?��<�
�{1�����G����x��C��{���y̆���/px��Uk����ث��z�77fgY9Դ{��E+�[a_��(��khL>��fu�V���_�o�0�������C?��G��4J���(M�⺂�Ʒ�Ko�{��gZ����"�:ܲ�Y]�Rg/��bUY��\�Y�?�T�_�����iuLN�Ǐ� W�ip��y�)i��gx������`؛<��}M�**BxԨ��F��o�85�5�N[[��O4��*�2�C���L%�ōWg����11>��ގG����/��~��^4&�RP�9~5"�Z��&��e�Eك'�^��m� �>P��_���9rD�>�м��7/djOˁʹ�NK��W��*}�n}
V߽��׎��S㣅�z�,��h�8fH��>bӠ?�S�O�&`��zj������\o����nę3g�G��׷�RjU���l?��.-��qr/���(� G
S�_X���\�Htl
X�Ǻ����"�=w����0�;{J�n
j���x�\���
�2@Ew��ġ�/.��X�.݋0�kL����e��7o�#��<؛[��M���N��?�ǫ��yvt\���3��|�"�8��L�|��t�@xż�)�޺'s�]]��<�
;����� �h�%��rMUa��+��+���=٭ ɦ��c�;::�F�M�]���?i���V>����B���t��	���vUҏS^X�������� z����Z��[����x<�Ss�t¿� ��>p�Õ�����q?d��S���u�+�؁��+l�'���j�s�ʖ���=��I7�
��z����{R��"���>�!2Pd���HYq�⏄c�N��Q�kş�RqD<��ӧ'�Tk�4���.EW�sZ���-�>�a�� �p@"�<�# ސ���޺���,Z[qG�*�/��O�/`��?x��5��i�c/Nn-�w�0b���~��@��!���q����3 �x�u׮]A=[]�.t$�=�3hb	fb���<,��v���|@1:*��+[�x�>�l�6�
��w���^��Gz�m}
�*��@�)�t;j��w���G�Ѩ�@w��$�$��ȥ#�������@E"~v�h��=�z|�+ׯQ�Sʒ����!��ޛ����Ii�b�yĞ���,���X�k����!W������N�gO��ѽ4B�6f��d�$SO�+T*���;֩=E��[vD���Z���L�Q"�!_�x�/�Y�w���Ɨ�w�i�Q���W�~�J��C19���Q^��ٱ&͉&e���@��o�!��ʔ��e��
"�YH;��H����@K�6�\�|Y~������	։��⢢�z��ކ=�������̟,�m_�]�7'E�;�R�>�*�/�Rw(k�x��߿�G�UVV�����
o�7-=[�0����py���c��F�>H��X���hZ���ʿC��'��MX_P�R����z25�g���J��"7,9@��G��AQ[[�����x�l�hS��]��J��o�@��!P�79Ih8u�'*8�CN�ih���)����p��C��4�v&Sl���=��8nȼZ���R��7&ዀ�!��=>�)�L��J�R�y~�O�T�o��t�џ�H�xI��y9���x/�`�V��3�!M���gv<��N��U�����
��m�U!�:����j�>W��9gqK��ʹ>��˅����q������\�m�ǰ������v�������C��)��+1�$�cw/�;9k��� ��~�냶�Gھ��{3P����)�oT7�U������Z���6h<�i��%���d��ǚ~�G8���+p
^�.��3�ߪ�b�������7�zh�=\�c��={�<P=Y~��Y��q�6��2R)���D��8��Zc��>^��#bu��}���fY�C^�����{q0BK���'�C���$��}xp]zW�.NN'oo�}�ҍw���P�����mjo�������6�����/�Ic3��;wd2��3=��L.���CP�W��;&�|��X�$Q�����w�Ը��k�b�v�̡�CN�3�Ni&��
�,D%އ�L��w%)�
e���S�^<�BQM-��I���ķ�뮿z�:ܽ|���e�d��Vel��FAN�5x3GS��@�����;$�zA:}���O֓��8�*�?E�ˍ�u����7�����!������� �޾�q�\#��d�����o�I�{^�x��rM���P/e�T�,jyb}Zc�!$��9���I�l��0ܼ{�[�������h9�ʁ��G!M��V�K#��ŉ�H:'G Y����6P�zB,�|%.Ж�\�?4�J�� Y���|p���1cu���ʢ�ᇅkך=��`@��g�AOOC�_5�rr6 ��({��m���)4o�l9m1�V,I8:j����E].��6�� ���C �A 8��P����e��W^�QS���L[|�~��=E��H	��φ1u�o�2W��C���x��x���X���D�� ��� `� �@�z�Kk��d�.2QQq
�Trko�w����_���(�V�D���~�F`��͇2�T�G�ȶ���}��.��̒��6M��O��=�Ѵ���e�%v�\���4����*��M�\6x��C���ܬ.�!��{f���oޘ%������XZ�G��L�G�b��q)<�+�NMM�US�k�{�Ň� T�-�<�GZMfϺ�p�OYA�~vͱ��o��Pm~}���{�+�z*,�/����{�/��9����\sBΝ���dne���Շ m��{-7wh���,*���܍����s���ۼ�4��Ws���o{|d����c�N=R�f˅#�\��jdd4���oP��[E����o�(�K�Y>�<��ĥWw�a�2��|��d=�իW�=���M �k߆��Vbk�E����/�o`9w'E���ΫL��[S!��n�0c�F�
M��@Ugx��v�k�?C�#�t4/��\�
$-�1��l�R��6�o��b)ؽ�V�#���ۚm������
b>�}��<
7��TZ��ԇ%r||�cbb���<y\-611��M}pjN�<���(w�s�$�P?�ɛ�*
�E��Z:�a�O_�r�l�:v<JK�1�`��
lnmM{�rϋ�ϫ���e�c�z�݋NQ��o�1�؛���e��w�#�;8:�hN}�<���9�8ٗ���<��o
2�	�|�W���D��Հ6���@ �c�����哓�.������D��gVev�(��{�\|V[���RS��-��e�үk;ӛb���&�/7g�`?0�� ��'��6aϽ��։�������Z˗/OŕS�򋻤|F�MFFF�mm7���3��3���Ibu�
�ۯ ��.f��͹��#Oߺ�����,]I[��`��5��n� ������].>y�~��T枟F⇂tJ|�6��P��.��+�k����k�^9r���{i]���~�"���\Ǔ���1�>����p��E[�43���Hi|�*����A�azS�LV�%W#�+ tJJ��_zS�'D�܊�E���r��bq�;w��ǽ߾}����R?P>>�1���a�.m���x"+3h�~�n!����ڵ���^�&��� ;��/�~�d�~x�(l"u�l���#���|�R�klhx|K����C?E��B�w��7e�����ޠc��M�4j:�i� ��� ��$5?   !���нշ��~�㛚0���P��~|>"��WH ����=����u�m_�`d������X�v�<W��-�~��/�&Bb;��Fl�g�w/�;�P����~�
���δ�����ڌ�/ޙ��?8���=�M޷�/)2KypS?��s�m	.��������U��oѪ-[��V���pD�}i�1PO½�U�S,���s��X�m�֏�@/�c���K1����F��y���Jv�x�[�-Փ��ӬT�7�����v��I�}l3��G#QV���}8Nh[�9D<���((h�(�L�-֪���oT�WO���_}�o�H� wT$Q���~~�j���"~u�qm�t�~�:�F�������;��6<�����lx�U��tYi_�@l��=�reAs j*��.ޟh^�{'��'��7���q��)[�bU	��(wۗ�5�4�nQ�8qJG��W�үg��A%&��+�������C�N|�+0�Q�_Ɓ�E���������mZ*����+=9[p�U��s�<��,8	k4�۷o�cr����zn������~�"0�݆=<��9Xm�c�TC�̓T;��ي`gh�l�v��IIe�o�ؾC�2�/kI�3sW��F�/RI꼴>���!���ǏV�0�&?z��p ����f7����b�
[��j&6������
�[5��1����?�5���QҔٵ��X�ʓl�l���{��K;����%0ln��r]�0lA�_�����g��aٌ�V�֋�t�������V��~�b���/Gb�0i1�xt�RUS[��~���ڬ�l��.Q�d ����2'�kP9+l6n܈�3דU��R�˿��u_�+&"ף�-�-[���5,@�N��(�޹>a�o��5;�൴�lc�L @�S�[N�:��8�EP�!,]�Y�*�@9�X}fh��~d^v�贝*�V�2DWY	fXX�_b�u �wC����]'�2�:qH�AL�(�3�ZP�xb�I�9��<�'�*��̅!�����dSC���]� t�=&&)CA�j�\]I�~6T�z�
X��(l? �x�9��8H�*y}W����}}{d��^M
	*"mx/$V������N5s��(���C?4y�oL�hvr��ց���Y:b�[�\��0$d��k���`�.�8w.���"�]���6�f#� ��򐈄���IH��g���+h[��r;%e�cmZ��%	!��X�@���9P���.����M�m��ނ����~4*<�-U��P�ņT�X�7��t�K���R�<��kc܌;����c�;��L�nX�U�	J4�dQ� eH��"9)93�"�JIr���$�Y@�9���'����ǳ�Qf����n�[]]Mـ��p�坽�0H�jۧ�=&��휁�#@
��Dn��Y[ZBq{�a�fg�w��δ&���}���a���H_��j xm���JJ��[+P���������/
�j��fh�b�U��+�*U��?v��6����+Xmym��?){�ȵ �4���F���9����U�!]R�m'T�Wl	_
&�+U��y���N|���=�9��>���f1�kN��`�����I��W/�g"�xh#c�w�H!��]��Nyyy��i{g�'x�i1 ���]oϡ^\?_%����U�N��`��j4��U���/'�:�������`Eݰ�ź!��w��gK~��y�
���b��U�����ͥh`��]��G�_�Y@��	�`�.e 5�����x�)�B�Af|�0T@�F�nA6����r�%��� :8}4a�0b �e 6|����2�I�9N��J��E_\�������|Ϯ$/J�z?�J�� ?�J�ؔ+ @ި
<�lL����뱿(a#m���[{��{���˲���v|Y�� V����Q���}o�e������ 0C�����ǏM
��d�z����g�GPكs��)����\���E�������|	�s�y{Պ]�[���Z{z�C�v>@D��eHp_mmmD�C�����w��6�MOW|/n�ng�#���y���t~��:���2������N�@R��Pel���k��iUxG�S<�q�R�2�nDd���>yBaT��:���}y��ki;�J��cכ믣��p$�S����F��Ҟ��iMM�Ʉ �9t�]iQ���:�/����uE"���*�F��0��9#��ϟ?aC@���8��g-U�'���g��:���n�I/b@� �3�:vI�[���|�UFc!lO&�����4B ��BqدJ'=���p<�1�齄�P��~�/R���{��6*q��!���
i&��%��LNN���%�7������k�G�P0�a�|��q��)P�9|������@W3���)A%j3�S�JP6��i�N��.��8�~��;^:�y^h��~��HB�C.X1�C�i�����2��� ��ځZXc�[bN�� ���).�������Tٽ� �F�JެP>���iH�����6g(������vnT�@6C��<*ג�3�E"��4�&��I�8��N���-J �rO[;rh��Zg����g�4���^}|#�q!�8\��^LB�����#�������˗�QB�'���z��Z++,�A��&�QS�_vP!+G�vg�7� B����Y�j���=z�Cv"M�VW�?"3���}6�<�/^�B	

B�70�)������(���1�����֚o���a!hX���@Y�77�T\z���M���P�1�40�	��KJbQQBX�� ������HZ���F.VQ=���.&	
</�êCR���`�=�&�}}|!�� ����|ow�9�n>��C�*4W ,���dj��&����� !�h߉������G�,L�z�v}�B�c������[)�䴰�_��a �C,,,J��-āW�+�S&�����g�߸���5�u��cx���;������
�K��q���
,�e�r�<(����.� �x=!/������~�CgExo�t�Tո. �a�0�	@�fg}�-�30R9S @�����d��)��Wƕ;�֝$um��i���W�~�������~���>�}�"d��e!�s´���yN�����e��C���$����d	`>��ɨ�Dc���}||�߁���)*I";�0�����L�"��zDRw�.G���@5@Zα������QUh���C��/�F����oW�TÎa��Xd$!�y%�H��7��6��\����G�3�s'`{Z�K	f��N�� ��}� �z��������\u_���@���<H�ˮ��㳧�����.��uN]���� D�L]خ�اpf{m���˰�"���a2hJ�ӯU숣�DY���*���,~��^XЁ`�mt���@гk����*(�OP�����yRԢ����A��'�؈���� 
��z��8���M� /��"��PƐ�l�wmmm
�hR����I)�Q:�6	DR���,m#�XwC�}Pﰋ��zK�T���sG4����5 +o:X��a{��u OJ�����G~�ػ�N�		u�·�'�В���	,G���|��
-��_ ��l�u�����P �@̀��@J�������\t2Q�@��KT\��I�b2�,�]e��wuYW��8I�!�I
��A1,,,%���7>�R��na�Y:�F�;X�E0�`T�t�
�oÛ(���;�Q��u++Y[[kf�ק�Q����y�+ѯ3Ka/bW�.gZ�S�Q�b���Y�����,L�'�n�;:����5�����_r���q����� (]J�7l���$Vo��>���y�����I1�޵vvj^؜t����Ot���#�� �!1����$$FH@X7����v��"���'`+� *-�G���F�p���Ā�-D�����6M1b�bG d���C<��M~"��b�:;;��v@�������O�āG755��O�
 t���г��wDxxZq��z-��x��ߪ}0���>,�t���Tom�Ѩ+q&M�$������9m g �O��i������;����`�C:����|
P���|"�,������ ��_�|�����ݎc=��;�מ��\ȫ��Qg)���r������+*C/���t7d[�f����>Ϥk�X��}� ���<����]:�΅Ċ
������ِ#�'��陙�1E��X��2�q\]u���=���a_��A4Z�L�F��sڀ�Nt�1���~���<z���Ψ��En�SC灷�X�~�n(
b)B༯7���:��&\:hY�br'��L��5�yp��7�8�d�m�YW`��ɴ�

bW�8�X�Zs���x������?�u*�ב�k��<��h�R3����[0٭�BAF��&lv���l��X��.�/����ܡ���˿�P�ttTo��;�@�Ng����qη��� ��� ]
<X޻��E	�_�B��+L�@��y�K��$����%�Z �28�3S]�_�*�m�;vjdh�))� .��׌<&�@���)�vD�=��_�5B�;B%�9���<�[������~yy��Q�0�.|�lO[]�\\K��\
�+��
P��a.ܵ�Z��{?�܆|�*|�
}d:溓T,�-�AA���<��OX��RIE��크`в��R���-�&��bو�l��"��V����C²xxdπ ̰l���%���f���o�����Jc�s��?c|X��������(��cA4�ar����J����M4�ml!i��mӐ§:�ٯu���H��f�='���cR���Z���.Ow��#��:�B;~�WS������f���z��nʒM2��4G7�����%n"E��yy�d�c�Q$��� �P��}��G���������y]\]��Ђ �:?�)*�8�r?a�X��<K��fWN������g����)�<�F��*ĻթBB"�pKO!��㙙��.���ʤ�e��l�i(خ�����A���ߨԹ��Լw�>i�g��C�=|�����@�{�uw�Q:'K<G��	�/� R^��F�Pc���<�y��Y+��p��3�;)��Ϥ ���3�a���H@D�	0u�:�%ȝ��,滉7ˡɍ���Ȱ���#�BK�Pp�Ѻ@� 8�<�<�Ȟ4�frE�L�{R��p�&�@ �^������n&���%�������yy��*�n�7w.8��\������6
�j����kddT�`�v��y���a@A�7�c�VVm�M�	���o��x���7�F���~� Sw��Y�%��ж7qm��y����o�r`r{�,\����%
�V����c��2�E6[O�[m�.����?p�YH��< X��pq���A:H��O��Z�es�TX?�r a��x���A-Aף�����l'�v�w.7x"""Rޛ�@����ʀ�p��n���M�_8�R���D[�4%���L?�@)�K�$bIm1�"=M�u{g^���J�&E(��L�&�l�c���*kȘ葟v���D��@��m��F�(�%xP�r?�㼿��x�/2�	#�^|��ׯ'�6��77�	Ύؼ�~�3�m�r������骓VO��)V֎��ʬ�����Ux�a�����߁�]�'�B6q��$[-()����S�������h��,�����^���<"��o�ʌ��vX�/%9��˱3@"���tD
�ɓ�F�n�TNB7t'��P��{ L��/%�Z��ߑ^�؂������] {#��^�{X��\�Fx΍��J��f;	c0��x ��?�w��ϟ�a2|��`����yҺ��84�9#C� �I��۷W���VQ��V;r�d0� �È��[c��޸��VUa�n3]���D��I������֖@/�\4�K؆�S(�6��*�x�RC^�����D1��Pɀ83b� sss�2/ ��HA�w"�L����$@
X�F�`%�K?Xa+�J�JX�C��q��DpssC�TVV�&NM�@{x�VPP|43�^2�E���\(߀j����x�a?P�0�7��W�8�q�}��Pn��Ʀp���lⱍ�? ?�`B�\o�	!�(LI���խs��%�}/;��Xܰ4���-������\�P��b�.�FTF&n�U�
�L/��^jr��6���<z(G�A<<�_�,z�%�.3J�I�P��N �:��Ba���m&҅�ZzzV$�%sP=%%��ɶ$���p�27��U��&��0Q��x��VW����B�J0�23�@TE�`{��zmw���#� ���HK�����^CJ�+&��@�wi�ۂ��iiJ�(��D^BX8�%��˙��@�7;�S��#]jZ65X Gz��w�%��2���cv�U��M���__�g��T���6�� L�?";P��` ,���G��*�i�Gڒ�����qqp?���aA�S�ɟ�
UI��XlV�Z
q��uH����g0˫o`@H/ANL��p��=�a��#(0R�ٰ�`��T@!y��L�r����|�e'�ԫof�%����,�92b<��8���1`_t��񪦦� ����^<��Z���g�����wO�k-tc�K6����LtW�q�~eK�H!x9�%w�����&Y��nOG��Ȉ��B�H��F�l�_H>�� /�+�P��Y�P2Y��E(�(:DA%��R ��Qd`߂1*� �A(��e�q��_R�!9��!}�~���0l�
�Ɇ��ۋX��.a߳I߽o ��ȭ��=��m��-S��W��[Q|(�N�Lr�����1�(K{��Z��u����4�AQ3yI�Q�j��w�H�"yS-0Z(P9ЅK�|[���A%�>����R�wkO~٣|y�l��g���Ծ���t�`Z/�cկ=��U���������W\a�<�qp��a�����Ty�ޱ��Ur����G�b^�2���ֹ��O���^	ȸR;�} �p�W�V򨯐G�
h9�wu���,�z�,p�#�+��lTu¹8��jj	&j~o��P02oi�^R�Z��չ7t)+�G���š��Ñf�:�QYu~���n�8�]3a.v�UGZ&���������k�@����*�x
}���@\��z^*_�����4*	QϠg�c�_R�X�L�85�϶,%�!P&���R8�'��u�ЫW�Ǚ�O�h�;s&?�3)�j��֫Wc����ǘ��n�_Y"٤�:�R���#�L�HY�����\T��cv`���
�:��<J�<���ϟ&���y�h����;@O�w�;���n*��JS�qF�P?ф��c5?��?J8:z�N�4b��u����N̨�JI5���G�X^e��˧񛚚�#a1�)�8VDv~h�'x���#r��<��H��NZH�pce�`�k��ꨓ�r� cɇ�L[������� 3d��y����������Ⱥ��6:!w�e?������\�+,�[��K/�~$j�pp�<�)��
@�2�cϨ�`"�Zb@��o�9jhl7�c��>�����e'� Q��������|����2ñd.@�h#�8����<~�D�Ƿ��V�5ӧ�����ob�=��{A�*��W��^�-��VTF��gs-�K@���ʩ����Hy�<�+ѝ ��e8�E6ڀ2�����N{h|zC�-��z��Pz� E-6���3b���gu�Nǰhuwz�٠)	Ơ��dm��������:j����Ð�I���U�|!�H�kR\QÔ���M'�I�d [h�P�.��"����vz��6�!:S�Xi_�N��2Ӗ��G�����[k�����ݲ���RR)�s��?W�OHX��[hτ8e����4�����r�dUWH�U�0\(l��������F�%ÖsM�x~Zz�.3�����5��"�$�5���f�\�8w�}�a'GXXY�['��ݬ.��ṈT:�[~�I����jc�qC��n�L��,���> `���[F*�TKIiEF�]��>^~��φOL�h���D���������*�2�[��7��W�5�X�K����_�N����5�f��<� l���]4�'�F�I�g�$:�4�����xԘI��]ӚuM�Q��/�a������L����������E�Dfٞ�A���堠`k` �~Nj
����^�ee�$��5�D�z4�(*!R� ws��Hw�o��C:�fGT R���������5�X4�Р��#����Q��i�j�q֥�++,��]��/�={6������rM�U�x��XD) �����LN���:�8�$[WW�"�㍬>�X*f�v�q�T�@��n�ϟ���Y�����Pє&B�nX�}kVm���XE+Go������X���V�p�邺��*-"�?Zi���y�J��d��+�x2�%��Y���X9��c ��ڣΆ��<�@��7h���\dV���7�(bN��lh_�g3����J���G�B)����J%�~�x��������sjD��+��&�c�B�ވ�$8X�^W�Cwi{xp$�֑g��`(���AQKS'#�O��^��yTuG#Ͱ�s�"���p-M�E/_�����5��ε'�YB�x>��C���|c^v��z����?)�f�!�!�o�jo@�y�0�8�bicx��e��\� U֬d�)Փ��<�P�֪�Jߒg֘kۤ�I˦�JϾ��Q��m��Y^̗�w�����/O�Dc�[��,�na��:,�C��GS����[��o��Y�;M�^��±�*�:����;c)u1_o.�1��������QQ���%Ml��/��-TU*�~.�K{n�p��ȑ�B��.��Å����,Z�u��5�.L�nIz~�h}����f�SD�u-pu���XO���ڗ�(_����pA���L�C�]l����LU+�"l��������ѓA�_���	"��#���%��2�2Ӟ�JA�t{آ��),aT/W�,�������;��
V�b��RB����Tq�F�s��{�޺.������?e�)��b�������t!�D�1P΍�*?�r�(J�,���g�Z�=�����ɺU��F�~.�p%>�J���`o��Ʈ?E�¤%�!6�@Yg�"�jx��խ�G�f���Xg���}����Q�������	�2��J���S5���~���U�%2���^�����ʛ�hS t��*�ۖ:��*��ٓ�1m{_=�\[:"��bar-��NH�����ď���"���D�d����s&ǌ�y�t���v�66H	����c��h`�m�y|�~y��ܬ�oV('A��>=���"{���ykc�fD�Lji�A�o4�c\���kn�Tт�4���M���4xs��rx�4r�Sc���Hz���!� ��]��L�C�O�^W����b��㛥O)#��Q���9ؑ��Q&�ӓ��s�bģ/��e���"ɬ�'c��m�%�a���l��wpbS��K@�&��N�gD�)�w�k���V�z�/z2l8��R��W�M.�ķ�����'	���@Ȟ��8�a3{�9��ۋ�M��S[��-�WKǵ��y�5�_���P�Zk���VYi�*��W?1f���!��*m��3�q1*_�\;�ؒEg���X�:7�q���/
sH���9ѷ�\��6V\�p��Vʪʓ}����ˏ5�i�NIW]m>�� |��� 'N����sԃ*�$N�<�=b�;nkg��x��1�<UuY�X�V����oDӏ�dwť�pڃ?Q���Z��*�4NB��=��Qǘ��4�Tš��@���4�}��H%S�l� �l��lO&���њ��	��'~s���Ri�|���C�w�37�$�C���Td\yu�_��L����$3YGL��C���� �&g>�.�����)��&��0>�(�⸓���V����XM�+�+��0���5�&����Vg>y��o��*�[k	`�=��_����W�N�,����j��O��CT\�����Mwl�=�(���%��>��I��s&&�v�I rJ��U�e�k��hT��?�(��;���n��\���6[G4���z� I��礖[��4,�[�;������<��F�&Bi�.Gww��[~����0\!�fUŃ�7v�T>2���Y}�i��G�:�}��=�P F_bT�1��+��}]�i���,:�C��]b�����c�^�^lޑ�/�.������G���l;���4xm�6��yF6�܂1�}�@��-ik)�%/ƍ�#���O��S!\��썔\�H�Z�D�wG��/ֺ�>P����Ko��"��v����z�R�ԸH��D����%R fx�x��6ְ[,����ۢGC�xA\<���[�at@A|�EEͨ���_S�@����e2���l�ӯ����;�;>��C8\��5s3� �R�!���ܜ������_���w��}�:����SL8������Ot�D ݗS�
�^��Tϰ�2�w
�9]����T;��,P�Lc����,�BV�2����I�q�իW�o+&����b�4ClR��$�"�?G҉)�{�r��{Y�o��r�������IӘ��:�Y����Ԋ����
��1��R�@,�G �tCW����Q���)��9'�e��U��F�IQ��Mܳi�wnX��P�����T7�O��؊4{��x����qn{K�J�^��y�Å45Ӯ��:]U��Eg�@'��W�e'�l��2X�i���-杙��ۂ������9���[;N�u��}�:mM�E�"�>Tz� �����PD"���S?Z]��IN�W9E7��{nn���'U�
=�i>�J�
�����2�J�&�9�'� �J��a\o��O���y5m0�&� ��7���7JJ�p|���8P=V��^z"'��п���g�`�`%�(w���%��W�/*�",�rqQ�?��z&�ag ��ͅ��k�q)'��h�µ�f�5һ��K23��u��%[������|+�5p�{Q����7d232��v�v�/���[��)/��l�잸*�βQ��31�;�@J��\�@�5���ϬՏ�5L\]v�Y��ز�9�B ���Y��7�61���D����ۭs#(���
9��S�.���.�;@�D� ^����w��=ȱ�:$w��V������R�=���hص�Z����IY� �h7-!&-�(M�(-�(M�-��&�v�/*Pb�Ґ��C�1��^/'m��Њ{Yn9�d�����LD�R��R���/���w�%���1l��2]��'Mt9��k��n;I73�2� ��/����S�\f�x��_�]�M�������ȕ�"�l�$LS����{i��ɋ"�s�;���Ҳ��m���`0����2c�(�,� `��9���-Շ���������|�+{�ό,���9���N9$㞸t-�n�,�P]�zvv���W�	f�I���蓵��)����Ӵut
�?['�yb��hh ��5ͬMcS?����͎���K>z�S4���˞z�X���p�<�w]� ��5N���/���)�8z(��1��V�b�7YY�Q�B%��ea
�uɯ�`h�	�]�CT_��~�� ��U��Ҧ^F㫘
��h�$}��V�o���Y&����=<ܒBl�h�s������jk�^X}��C��_cA0Q�gK��{���iOZ�@���}��aɖ9�^\�p�Wc�P���QVV��	->[��(�|�gB�#����	�Og�����b7�ucгL�+�9��}�)�T<��uO�bN�sB��Xl�ᯒ��/o����1%�m!��
��;��[ȸ⧶�7]51�on=ۘ����,�Jc䳛Ӭ2����z�vR'6�34�;٘ +߂?5�h�K>n)�I���U�"�ۡ������<Hy$��]�?�b�*�V��/�Ԇ�G���4���#��/�đM���$x��x� 2+e)Dqc� `�j�� e� i��o����럞dm�g��Txm5�Y8C;�/��
�fs�Ԧ���N3]v����+�|V�К��s�<1��[W)�rv|ثG�ir��<1��~?��q���z ������'&��K�H��iӎ	tN�<���C�NJ����B�#���qx�l�:���W����Qvz��}��lE�~x7��@��d����T9�R'v��5�x�ڼ��1b��sҳ{���0�SA;��ʺ�Y���o9���0�W���ӷ���w��7�-滖{e��%&�� X��"�;���<���p�g�H�v�H?�->����.�o�ɾ��xG��RrTǫ�R��`K��8��u�YI�)F�9�ff���v��������q��,�ʴ�N�D��R�qW�y���>���r;������__H3����:V��4�ބ�~���6I�dO�-2$M�����RN��.���B�U����w����'ؓ�6���Q����zZx�w!vn�*����s4�v����fD]`���ä�s��%$o��zqf�?�o�`t�n��f�̅�5�U�.H����!=5!G�"6]g�"������o������^h�{z{~T��d�����T���l��3"�/����,�#�Wz:�Cf���+ր��k�1���/�n�,,�3*�s�ڗsm�--!���U�<R�EM��Yg3��Ɲ�Vwu�\/�#��/��B�trr�'dǮ�m�/�.R1�F�b�n^,������4�v�<����8�#��x���c-�d��k�4?\ln�Fk�q���|?��{���|�������P[�2�d�s�����Ǹ�_vu��`|%��`�b|IK9�>��`̵�k�*��TM��?.��XЇ��"���±O_T\+�c=�H:�N8���o�zSN�����\e&#�����.��(oc.C�-FT!�[k�D�Q�Cu� S�>M.6�/�Nj	*)�c�y+�fљ%)+�MW�bW�f'�'Q�S5H~0�	'm�j����=��[S������l�K���mOr��ƬV�nJ�vdA$ZH���@G���T=.k�F�K\�ƻ�d%}gV�MԖ���S:Cm5�
��n=�[��9�t�SNM�gнYgf��ga:d;B�;��%���b�=,:f��T��x��1i���/�LFE��_��~������?�}`����0 ��3�v���Ng_���ם�y�ʜ�dZ��cF�r��bP�@�����@�0��~0�g�c/���h�r�̌�t;V|�o�U�uq������A�v�zc�u�4%�P�!G#��gg��d֫��"Ͱ��g
!؉�li������+���60�k�3���gy����y��`����9|�C� z,-W���W���H�I/��`;��?:n=�3�e�h�1B��z���`NY{��6�9 *��d �`�֖� �Ǜ�h�ء_]�`vL��g)��SVL������3P�.��}
�ea�A��\�j����n��`��k�J.<m�	�6������Ϩ�؃����������'{i`�����өy����;��O��k���8�s�f��8��B�$`/[� �澜C��h��+\ݮ�y�N�Rp|�����xjwt+p���W8y��O]�S_����Qv^ǣă@���<�1sU���ypg?��Nޚ��$�6{���v�9�����u�F���xI��hifZ�]dpP�n���i�1�R��G=�:N[,���β�q�����a+绛kg���Lk����<w���<cc8[��;f��g�v�8Y�.,��(&*���j�5�!�D5J�l�_�~���﹟
㓀?.���3Łu+>L��=qJ�
Ӳ�޻�?e�QL�+��a-��әҢ烵Y���v}�4�`��F'J��K�S��*����8?O��.�������2k��̺P�D̔�P~qqZ�EUb�"�I-)^YzN9�[4�Wb(Ki¼i��}����=TVt
��b�0Q��,�?��hc��\85��c�J��M�*uވ��"��h����^����� ��#ƿ�߭��0yasA?4�"��y��Lp�1�t��|�M7@.������g��#�fL��ڴV�5��
&�/6����� ����9�՞),D��#`K~nq<��N�����=�Q��r��3�cH� ��v����f�E��0����3�e��<�nK�r���|CߤO��_)7^wI�j�T޷wޑfπ	,�9���VPP�@���]W0:QIOwBE5�t�ǯg�,��?�d������Ga�����8���������j6ݸ' !l�M�'V��J'(6z#;O i���δ���q�̀��j�P���R-g��b6)nҐ�KC(�e{Պ�7��������i���L�6K��y������)�g��f�����#'̵Fa��q��@���-�P�����a���q��ȇ���u����8�T(�f4�d�h����R�vܒ	�Ɓ'}}�v���lAR�F8K�D,���ރ EuN&�4�� ��72YN�ӳ��֜�e�)+��ĝ���l��7���1�)(�7��V�}����,jy�1{����TT˂����W3�-��9TT9��D
A憘!^c�Q]����2�`RI�����F�8�s���L��x�.��";Y�;O��X�Q����t��v���'�J3�b��ơG$�ZE ���p��E����ƫ
�pٝŦ�&�z��kٚ���{3�ן{�:��n�j0<8r��}R��K�n�4�P/�Z ��yx8�D6#����3��+d��T=d�G�2���^c����8�P�u�E l+A���z�Ų5}�C]��ʋ������C=��oő]�����2���\��xЉ�f����Mb>N��P�������e�C^�|��qB�I��StH�9_��\A:.�kR��&s��0��؀���Fk+��9"ɺ =Ҽȗ�h[iy�����je_i��l�����F{�+FH�*�9��^�iŬɎA+��$�h:x'��f++��U?�v���Ii��������I���Ur"/�r��zfM'�IM4%���e��jYҷ�e�7��q%O�Ctן���%.pCr��u��>�B�� &	�T�G��P�b�iv�����\A,�l�Ȩe�n���1o��}6�$��t8[�e����{Ϣ����Izr�\/2�"�3ѷ`�'����Zv�;{����7����W+��%	>��?7Lr�X�!V��g�.k����&Cfe�v��ۮMuK\�����Uq�������?���x�B�� a�?1�T�OL!�Uo?���MTU�lA��Y0�`)ջ��ie�o�!SV���kb�H)��Qs�D����ª���kzm�_z$+I#և��W"{����� �e<3��8z�(\�:FM����Q5fvr�����QK�tA׮ )��$�c'a㙾������B��������Ѱ���M&���{|L��I N*��n��Te��@��ʄ|\��rj�y�	��;�<�]�Q�1���ǽ��JpWۻW�$NĻ�.�,��hx��Ӑhb��HGJU�*�Kkp����g\���]8�I�"��������t����y�i�ػ�J�<��y�&�!�p�*+��BF�[a�v�xz�6���/i*��Tz_�f�307�����P'�V��63�ʳy��S�Oߓ��"����#���2���kpv�3<���3�:T�x�v�JџM/����A?À`�q#�E ��T���kjY�z������jI�t�*�>\d��
I ���o�3x��_]��B]j�-��УZͽ��ٹ���,�R���]�f�=?^�`���<���ߨ̓?e)��R�''����,��u�|���
f��.;�}�_���J�VQ
��yrFT� T���͗�X_<ͶQ�oRà*���W*�w������x
�s�&��	g�M��t����;7�!�R�g1c��n����M�F�����׾&N }r���@��i
�Z�x��N{C�'1`���Ϧ�95��Hym��<p�ј��5�/>�l�R�0�3c�)ݨ�Ȍ�<�� �`�����4 nIea�?�1`VEX�ɴKL�b=�]���t{RԴ�=�r�7��V��/�#��a�?���c�`4�����ܽ8ͦ-̶U_iS��2�&�geLo�n�g��Ee�����9�0�J�&�'B{��=y���Zf
��2q@T[�Z���lR�j���;�k�ǻ�dߗ|#s)�f���ꆪ���O'�m~��Ɠ��.k�jO�)�:��������k
�P�'�G�<V�ÿ� g���y��S��SN-SK��-�@��uD�W���5Ͷ�?��FW�r�Z��� A��c�6��H�T��Mʯ�D��a������͸���)��IQv�EH�ՙ�TpZv�����[�!��7�)O��
O��ʯ��x��u־�T���`���o&����������]�b�ȵ,V��Afw�o�!�⾮W��.]�
�aQ}���(S�EQ��) 5 � �����B�մ���

��?F;�:)y�Z�֮I�Ƽ{����&�X��ĩ� 7>�Y"�k���9L |�c�	ƣ	&�)�Ƞn�������6���n�Ɇ� ��ȴy�X��V�@�Gk5�)�L�¦7ަM}�c^�b�K�4�m��)�[���B�z�TG�Z�о65-�01�����Hi&��h�a�iB��G������Ezp98r����/9t��VL�U��������*D�Дb�9��7��=��69D�g��_��)�̀-��:n�!I���B�Cj<�p���s0#��9�.
��/7�L�}��Q�M�*�G�c1�]&(�_'*����-��{NV�o�@i�QyPN��o$��ef15����ӫ�M�k�
����s�Kmg��L����!S�4����"%�ͧ$!,I�
�I����Db�ru��=���g�w@z^0]�� J����>�c�B�+�e>?ʯqFw���[�ϖ��fژ=�� >-�G��S�W��oɓ&����K�`�NX�N���zRP���9�c�J���\���>R���;-Ast����wx('��Y�;��v��}�0A�s�ӎ=�r�FJ�S1�QO�br(<�S1��ӤR3����X�[��F�[�H�X��7�r'���n��`��.iSL���r
3%���w����	u!C��m��ÿ(4������pz��0u���gJ�F����R*�M��M�x��yk�j
q�݊��h�Ĩ�qV�����^�?Z�>��5��":��,I�2�۫�w�ϾT��A'�)H <X@�%���l/۴a,�h"l�VUt�ٰ�c:�j���5�~攐�����8>��[���V���	9�W��_C�x}lz�Z�8� /��o�U5����"���j�*��	��9�����6�j3�u���UC�mZ�B�3�?�V�9�=FwH�sڋ	��`Z]����ȣ��ڱ<�lt����i_OO+��"uo!��.��Ƀm� �K8#k��f;�{s�|j}pl�sX�JOM@��v}�
7�2�������K��c�[5�)�򌧜�]�������S!~�Ie����#8�p�sUaLLL;XY�n�x�0dYC��
uo����;T�d�m��l���k3�CL�5�����Z)���.�o�k� �T/����m���2���o��]�UqUa��T(��{.KAUV�<h)�l��E9�R�{L�:O~x����A��Y���,z�Q��[As,���O�o�
1�Ƕr���W����v�>pq>���I^���uLP�}��ѵ��������[��_��|b<9�Ҹ~bSyB����t��VF�`������,��T`���r�.��igx�4I�}�SA"���$�rg�� ��yUL����7�v�M� �����S��ՅŮ��%�D��Vc7�nKS�l:�jLCD��p�t�
�hpX�J~��Ì��C����<oG���u��A��/j��'
*|��L�E�.F�JA6��f�*�.FG�~=KA����M-�L�{�h�}��/�y'��� w��|N~ /�+ϱ��	�vn�M��	��9W��mzӴR;�U�Pf�lLJf��n���H�IT�f��0c�bBb��>f)�kS�c���,�w.�U��	9�B�:�>Z��w#̀@���b�q�E�M�J]�c��l��gչ߻�[��t�xٌx�{�M<�UK(т��1���8�2��G�$�:�Zd��Iz��T�������,�#��U*+=���)�j(���]�LH�o9�0�̰��Վb���� ��A|��A��}l�*�V@ ~w-[,��tFִ?3���U�lz�����:��:������R����$����D>���zN6A]�
�^�QIЇ(Ed�Y�aRS�i���7u�ƙ�5\\Bb��?kve<�Ol#�X&�10հ���@!{�=A߬����}>�m!��H�y8}�<�G�a���	-���熛I�^�1M�-)h��-�3�-��g�5�5�O|I#)w;l�� ��?u<��,��~Ӛno��E��]���� n�g�#�WI��������Ku�
���\Ӂ��I��i�P$I��뤠��;@,���8-ױ��iJ�v�Y..n?�:��?6lo�4�e\�=�hͭӾk�'�&JU�����6����!/�q��p���,�NG)"�<��h��������#�����jfh��Jf�l*�[!|A��� �*�wS&��>����I�x���tg���f�k��w�[h !��:��O�^�9-�$7J6�O��v�E}�Bd��hB/ƇormR�F�&9�G�<c:�ri�3p}/f�4#�� i�*j]��YX}CC�Dٳ찲L�����Z ��ʽ��Z>o}�Z���orr�i�!i��\��ߘNмD������+-�: v/�m�H��!A� �X:�{�]{QF��BO���-�u����'�U����7�RVF�PC<�o��k� ��ş����Wk���D%V�2�{ Bd�I\s��R�F(�Ó[��� ����7�L�}�nq�y<|�i(�W�i��������g\�����b�+��>u�����苫r̓{�ȵp��&��� [^f��S����:��$2��F3�r攺�����}7�R��1�G�����y���������je���a��#�8(M[dv>��s���*���1���ǘ�vw�z�L��ti	�x4*�[XNc�u3�M�h�Q�f����	��;���%�o�g+Emi��H��|���J��H��p���M8���a�G�k�C�G!
�����������~���Ht{P#����V�|F���䯑�R�|��[&����%�Y�;	6��@+X	LI�� �_�c� ��j�q�qFKrP��_���g��Y�������/M�ca'K}�����u|��u63������ݯҋ����^o~v�"{p��w�ɞ`b�$���	��Y�lyt�L�Y�d=[z#]X0"�>�S(;n���a+Ol˪��=oAp?an���Wt�+���q=�b;�Э���TT8KI���Ǳ@���3v�qU�)4��o��n�c� ;��-�\�j�\��D�8}<��d_ܴEURP��\JW{�4���U��=�9_2�RK�@���������j�����ɦ���,=m#�����m��Q �3�w5�o����<q�R����Y�.�L����*v,�����h%R�a���6����Z�E7#X�mZ���.��p��Ն<�4�ns��N�!�0�M�`Z��0^�0���M�r� Q��n�������������ox��D��R�z�B��l�'�z�8�.��ND���z`{[�hoYd��
�1�=���/��:���M��R����(
��BM�D�$�%�d�5M�B�ވ�gYBeI�d�ٲ���;������3�y{�^�ܳ<��{_��)�y*B�f���K��������F�l���IIIFj�ed��߱��ח����Htkcr���X�^=�e��.|��� ϐ��e�ofX��Lz+��x�s�b݂gF�%��;<�ڵ��*׮��H���PMM�!��(J��Wod����0����o��&k�^9�?���Pc0��{<�\g�,��W��}�Ҫy�c��j�ո	�lƑZ]�u��n��Ƙҋ������>>uib�1���� |���h.ޯ���y�V�鄔#�I��r�u�᳻4D�t�T]k3;���������Θ1���v���ҥ|k������Y���u鴤۠4n���b���%����}�z�#՚����B���� [�/u�.&&&Fmd��}nӍ�T��d�l�k��4>Z�޲�%:�bb^$'>s�v~����������T�.��/�n���ԥkH�~�������d�	6�#_i-j�di�L�~���9�PR���࣫C-�&3�dŗ��Ō����Y��1���.���\�LS?�k��K٩<�N��h��z�7�Y�h��o��M\j|m"��%7��vJğ���y��Y�ً�n�)2�;��������"^7�:������g<�F�q�)~���p&�"��'�Z\��<g�6��1�l�����J9S�n�����W6�j�Ƣ�j4�_87X�LD+���tkLOO4ۅ0��y=�Z��s���t:`�m:��t||���=I�Ul���.�����_��s����ӓ�����o���ï��ދ���w0G@�.���{L��q���W�D(��=�s���/���=���];~6��N��/w��U,�n�j�d`⯕��.�Q���r�{zD�����9Y�-vx��z6 �%~aҚ��9��RJ�� _0��|+��c��]Z1#�w����5L�Xv=zd���B���k��,�v�P�Ն���v��5�w,;l7����*7#������q�y[���=����[��ol��X�����F!�4���*�OT�;����2��ܻـɩ*ߎ~�H}ˋ�]�@\J�<��·� Y��J��wzys�ߟ�ΎU�d�<rƦ�V|��]�j���dq��i�l���u#:�����M�ͫVX�V��Nc��_�����*/`��}Q~#X}��3Y��f�l n�����w]^4�o,;�`�_��6)8�:����@�L]uL�^���/Y0�J�~����y�o�bzƇ\/>��� ����=Lo��!.�=&�-�����+拄{��Wy���H�o^�`�ӿw�8~�g���6�:���/���Zt�*>�\����*�\���:rݰe�|����c�E2�j�.	H������ᙙ�/�}g�9�M�/�t��L��,�En�2���;�&!�c�3m��@�v�O��y�s\�t2�o�a�K�2no��-g~u>RNf^�������m��y~hP��������
5^�������%���/�S�%�r��mL28��-�_S�-}`5���l��\��sms���#w,��V�[V&B��Kt�Z'd�c��@QF�Pѡ���?d:�?R���Qxd>O,+��k�[L��x�8���,y�n,�h�i�!����~�����ꐐ�f�a9�n�yќ���,K6Ez���ױ[ ���
�\�xHm�Ȼ%�

���q���vC-�w�`�9�������(��)�k�~�L��|c�{g����?�׌��Ͳ�O�j/�tx�����=T�	����F-ZC�9ӆ�>���Ek��ۜ3���-�r��\߇aןM��\G��au�G�-�7��	d�ճ�ۏ#ڿ�i`zd��ЏG�wx��άʙ�'& 	��#�k=�dr<ȱܠL[�*=ykD�,�@҈۬�����~Y)W����.r�,�낶�t��8;���ZɆ�S��^[!7�'��?7ƒ��a�V�.�g����������ٺ�+mQ�v?�8�{�;��}�ï����*�X����W+3�W�i�l`z�L�S�%wy���������7:\F�rOrΙ�Y�cY]�A��%�IF3�2�i���<#/h���������Zﶁ<.�o�s�jD���SAY1;��s��f&�����"8 �&�*�8�rGw���Rg��m>=���]�-�-O]�9�x�i�SwG��ɱ��(h��p��Z��%�xf�~Y����_ڜ�·�bW|��?�<=)��]�Z[��M�,�"�BdɫrEO��aW�>�c�� ���Y�_�.��:J>��z�
g�9����tk|�my`|���\c����-��ba�M
W(ᱶr�cꔹ�7���S4��*� ��E�N1ky������O��>������0�^S��yӛ�Lҋ"_@�zmj��D����j���_[�V&���}}�.ݬ e�쥜����?��h$.��8��*���:A��;G�\�g���K1��*�U�w�o��f,~����Cf�92�-o��;�q��R���(��e{�E#�k��*�ҕN*]��t���9���,��x���&<=/O���f�]��,;�t�jHB��G��4�>m��O��"���HZ�,�]�Ƚ���v<�5##���Tt	�e�6;5^g��\��r���x���M,9�ԝ?1�w���B��H���RR܍��Xa��8�����������{m�m}`xFZ�G]�u��,�Vqu�20)�a��fYܛ��^��,���h��{F���6(���Q��rؙgZ���DH̓C�a�]�R�t˽��Ѿ߮�վ�O��E=�y�2��1���1*��:�#%�����6E=1(�$���~��ik��3�|�@� ZO��/�[�9����չ��rS)cm�J��M������i	�1j���"����of����
���14-�Ѽ����8v&?Sݚ�n�%<�\%X:@�r��X�%K ��m~Y���q�wtW����d�/p	K�i�c�4~JX]�>(d�ޝ�5�~W(L3���9�X�dĉ-��ϲ-��:9'u��p?X���Af�
I�'I�'ܷ}��(��`Luy� ��d��a���.���~4[���aE<|������I�vF�L6�:K�9��'�@�G����/8?�d��V�&S�Y��,	K��@#�4�0'��k���u�lw�	�[��}ť.s��GF�x!��S)t	;SL�V����)3�i���g���OoD�/hL'�F�p�xk~�A̯zg"����z��3*Jp
}z)��Ѣp4|�ڋK�w��S��1؜E�����`j0k��$scQ���@i�S� [y�s�1����5Y��|����(��H@����J����g�r���鐇`�bo�Q��5G���p^c�(����h� 7!�E�022�oL�����S�?5�S½�k|���i��`	��;._Xf�WVZ����+��GWY��6�B��ɓ�z������i�o����x�8�/ϼ9�}zbH����г��@�x�1Hr*2/���O��he�X�$�� �ffJ�'����h-�(���VE_���"��^É�1#S�*����>���6Z�:�.�,gn�o�g�u�(�Ýa<x���d'��lAJa:?���%���j���_ @�+�z���'�W���gn��N�(v��$��i�O��W��9���Uֱ��׵�LRz�L�SR�����u	T�-�5�w���I-�9SLФ&��l��`��_rI�4��+K�y:w����K�kρ`\i����P���p�f۹k��:��i3���"��[���W\��H$�3^Rv�Ȗ�"����&[���V��n5�
����P����m�	f,a݈!sƟ'�`���Igf<���$�"(���{m���7���[�(�4��_�c�Hd2rt��j���6����S;� ��D�H���G�=8!�+�!���)֜��Wn���J�cĥ�<���̕��x�^UUq�^� xD��cl�����r��>�����[�)�;Z�}�m5l��x��]�:\m����|���z���H8�OE��������O��n	�~m���	r7�E��5�>&Wc�L���JR�n��rc�W���u��6�/6��С��ڨ�3�;@���#��2Ĉ�A�J�I�ٶ�6���aT�UU#����r�>�sދ�	��vt�~UQ�v�A��?���Ul�qLi��6h��[�Hv('���%�_A%	��Vy�:!��[� qT��ы�E��8�%XE8 �E�;���Ȅ�Waҿδ��;��cvf&�_�H����K����;R���V�6y�NOѵ�Zl��{�Nl@��u"ٸ��U��샲;��o��hGx7NRU��V�P�HB�]��Q��Z/��Rp��Ԏ���{r�W��㾭���Ub�B&���H�!�����_��Fw���t��!��l�)�+�rg��R�����)ہ<</�p�ۅ���o��*�L_t<���"nU���#I���w��� �(� l�����@_�~Y�y����Zp���Lk�S��Q]>���=�8��~�צ�U��ik{@&:��x�h��'�����=Z.E!�~Հ��3�[	��x� �$��0��e{����P��ޏ��'�g�5R{΢��V����8�
�=0�E�:u��X{$Q�b�^���S�!a�t���n9�k��s8�NP��lB�p"�3� 8�̔�llB��B�h_'��IZ�+�dZ�a�NB���-��h��.nt����{�����"�:�Y%�8���0�]`�/���5������{�?��)W��g�h�b�ȕ���@�h���p�u� qm�W�Q�b���;�	&�?��J1�P�+5�YMU���5���OJ�m��Tay���������m��<M{oJ^?��$��t�%�@:ݛ.eG�|u�CT[8T-��9������<�.���T~tو�3Me��:�8��G���i��`����w�m��٠�>A_����R	W���&8��Q�eM�� ��γ�u����U@9��u�ƛ_�hf�*#�����h<�	@%�*!7��-�d=������T��?�Q�6����n��qzfB\��W��D�N��"�}ޱT$���s����bBP�UK �����.35�`�dީr��w��h2����EP�?�_ߘ�W!�,�5!B9l�ξ둹��E��9�9_z�l��@}���y�C*3��Ӆ�ڇ�/�L��#]����[�NAݺڢr�=�����7�;��`��Rs=;�H�4� k�z�E�U���x&a�G4�j{~�5�==���J��?	�����q�P��\ߦs~��v�C�&%&�'�~n�*�C��S*k��uN�[iЊ���AO4����H7`cERCُ��It����o���j�����q��\��G��FiA�
��p��({�0�l�ך��@�d9�j�
fH���]b�l˥48�;�]Q�u�ŏjG�ȷ�ŏ,;?�$|湚?�y)�A� �|P���"_�7�Wy��W�@{�[1=7=���+�B_�k�l/ ��Ϳ�*<uҪ�#}��Z����R�x)��E�yL,�Dx��g #(V��h�������T����6XHc�~�S��	@j�:,���/J����E?;Ĝ��;>}S�:ؔ��+�
F��rJ��S����k�i�����m�W�_��lGF1]����o	�.eR��">�������]���� y}H�
Ņt��wKx���{�Hl��Z^�K�I�S��i����*�L��@�5�ހcV.8�&>���E���;���ہ ���*T5�	�-z�`l���Q\N�7�n�Lz�����@����,L��Y]�:M_��2�y&�b�a�b�ؤ*7��${6��X!�^��\�H�����"\+:���m��f�n�sl�L]��F�� 1-?֋��xl7A���ȳi����J^5�� ����$��U$C?�r�w�oL" ��Vޑ�C�m�Q���t��_���`��YH�AM���H['ʥ��lX&��x���Rrc�|��@�Q�m�j_I��أY���B�= ��+�w����7����e��}}�~U���F���4���l�4�@z,̰�g����H�17�R�_��U�Y],�9k�Fi���JΎ(�^����#\뎊�B&U*@�M��O��[��̄#�*|����ͱ�1f)$�}8K�J��U~�5¡1�o��^���;��;�@����_r36��ƬAA��l�e�2,1�K	2���C�%LuY�7Z� �]J(��d%ˑ�PRV���}5>�"dJ��"<#H����WD����b�W�M�&vkm�g�+�L�2�T-;��5q&���N��D3��vg�T����aP����bc���0_oU�cD��j��D�qe�v�N�2���n��/���V3�HG�����f]�v虜�,2R�g�!�'@KE/�?Z�B ،�<�&�ylT�i�t9�=�it�cEe�(�ȭ�$ mF��졄P�[5�gF�a'�Z�q��Y�ϳ�5�o_��ӥ0}�Ɂ\�1��, Zb� �dL������*�4drCqZ��w�[?"�����.���j��'ٔ�h4�����Gp�ȳ��[t���'>�g�����魮A�L����x��=�҂�1z�ǳ��{7�� T�,D$md;/2?�]��w�ژ9D�����觗��l�gtt�x������-�>'((�$���n$�ð�"�(�]���{��0߻ʂ������[�g6e���ת��&T��Q��`�8�[e	�%,�+��񾺎�hu����Hv/qP�£�|�
�C�M%��[��.���^6������Ծ������QA�!8`���?P�ʑҲ��y�Unʙ6/-/�(w��$K��G3�٨���w�v��I̔MV$ e�0�H'%�L��s!�$���%ؓP"MsZ�^�ƨ�\�G��1�"���R��BUI�V����XO%��r!�4�lݿ	'L�����_���/���d%<ܞo=8�y�+���D���񮝩�+L������Q�ǳ7��`���v{�`S�x8K����I��@��4@�r�k*�D>��|KX�fV]p?���6(� V�T�w��M�CI&� �Yv�-�,����i�.�<XS+�Q�* j�D�8�G6[�����L�"~�pZ�`f��{RSf�+N|`Ү�W߀O�(�%)k��[ۃg�6�\gF�@/B��̞n�,!|�6�����%ȱ?���Q[k���i�T���������>����� Ly�X����"�^��R���k\{ .���� ɝ4�B��&>���}⸼�/4v�DF�����QZ�5`�r�� �#�;e,�� 
��'jD֗�O��Db���*X!{�hL��bv��X�RŹB~�B��2?񐔼-1O�'Yf�B{������0�;g0q���wl`r��D��;�l?�b���Ͷ�����,vV��9��\<��r��-��R��د�qߩP��j���O���>�/�1�,Ј�M�&� )�)�ǧ���ԏ��4���j���h,P�O;�X�wy	Pu$Yu��ʿ�Q����=;F��WWO\O��y?���v�$ڦ:226V7��F�Ȁ�l7�fLd"�r�H�ҽw���m���-�6���{ ,��jv$1\�FZ���
`��Ϳ�sIX	*�8��s�˖�N0��ig�D�ς����\MT ]�nÚ�x��v�anO�����ݿ�x�>�T�X1�@��'\_2��\tצ-���Hd���h����喽_^��Lu�����͚���0\J��~�9���7��&�:g��S���3fgj|�fNA�]/��q��{�'lv,t*V&X���߿�hI�w�_��la�U�����#��6��${�f4�&dZZ	�'`�N����1l�����"�J��!E�|�5��FFۑ��'�`ɀ��Z���4jPfo����]�g����������b�5��B��5b����[R'GM�x���R����&�0�x.���h¼U�?K��^�>�E��އHzh�#_�Ep}��p�6�}�S��I�N���߭�&�������8�L��uI�a�5M��~5��9.$W�w�-�Z�t�(���4P��·���' #mu~� ��s�]�$/.Kފ���W��qS������Y1�!�8��W�v�z׀j.y�y��W�g� �n�i��Ͳ���V�x��=3{�G�ǰEZ��0��l0�jȰ2�Նr��2R_=R��������@c���f���ysm3*;�w�災%�on��*\nPF�^��]��O�" S!#��8�h���:w�bx�
i�_��]N��	��/yksrb�%�	����q��
~{Q����Q���ݐAmX�a��?~v�`�L��wF Q�}��A£���;��g��6��A�Y%��e�p�Q����k;�$a0ʢ:01��`}���b�ױ��Ó��~��@���K�$Vs���>8X��M�X�&ڋ�LOx��ȝ�O%3c�}�-��I@�S�bWFt"(�e{o"������LKpYٟt�X��T��ǋ�~�[�ل|����+����3����U��"����>V��G�K6�)H��h�q#��8���l��ɩ���*�}:�l�dD[v~f�hm�au�{�vG7���dS�b�׷N���k�P�xı��r�tjD���>��G@���˷B�^��2�F�Ǔx����+����� 7�7V�٫f�y�@�h��/!�8�;Q�}��?/�X&�6���>߬��Q�#h{���>�wWߊ7a��ގ�rTL�@@}`����4Ǔ��I��:v�=�n^@*K��*!`̸���+xӪ����b\�M��	���x�>rc����F �#E�6:	vg��DLKV* ����+:W��vI!ԏ��kWi�o9�C0<���{��BB;o�:��O&C��9�홹|��k���զ7�3��b�V4g�	�v0�(�j��OQ�ݡt�+1t3��$D����h���� ��8��)�tVhcϥK�?ho���≶nUU�p"�F��k,	+q�n�z��:��{���mb���5�f����q�Ӡ��h���������Z�����,�h��%#���l���!_/p~_b��j}�Q9ܮ����s���)�� �u����י�rX���)�����ҟ�?J�Y��0)����<3理u�I�^ml���y��^��n���'ˎ�6�3��8=��P	_�f�XrR0��$�}"%k1��42ĕ�n�	w��dA]�Jc�_�P*��3�� x����'G�8�x
�}rrC����Vt%e�
a8�r�i7�`��+�-Y��(©49:�gK�ݐ�,Xn�8���R^&�lQ��.c�<�7l�28�6�C�O���| 4
��������;��
������4)��:DM6�n��z)�A>� �#bv:��ΚQA���eE�!ޗ�AK��$�����i��B����eSު��''>����e�Lj%�?�A���:���Ew��/���Q���]����� �<rɖ&�& x��ߚ���b�;����Xa��ܛ%
sB=�,:���ju|� ��Y7�:��-�9\��#�2Y�J�o�@��$kT�����������y���7�$~�jH���&��F4�_v%`����I��`JFת��T-�਄�9I҅����!��'�m���ī�)(y4@��pV��vk����/U.��;��7��-L�s������p���C�E�W��Ԑ|��F��QDF���"�����H"�w؛�M���Xh��Q�/�?���e�t��8�F,h�����"7c2��"Kִɡ@=;����� ���@��t�4�mw=�r��1�V���d\���c$��L���dg	p��_?Y1,s4w��7ٍ�\���g�Bo�-5c�nr��΃(��i�fɺ��WTdj;��L���*����ȳ�+�3	&d�SOȷb��4�}B�j!;�]ƨd���e�,�y�2Nd3S��.�9��_�:�ʖcg�-�W�{�#6�3!6���ur3Çѷ��y���FJ�`͗k+�i��z�x(9��qW72V�n.J�}�1�#�&������g����1�p��
�i��H��¡\~ҵ'^S9#/�Ӝܯ�8���Oӿ���ʳ0w�Tl���Ti���������w-�¼����MR*w��H���y��Po���V�&�^�kK!��j�h��-���&�^��N����k��[g�E���sPb)��,�!^���A�O%������g)������!%�󀾴�����VPk�?_���I֖˹m,))i�>��,�טq״I����;���+�-U�;�OC=�t���|�O�z,�Aޓ�3�$�_��kW���S�]f��?�Ĉ�(൏�����8�\��bdo4vC��H��f���7��gR��o���7$�O��T�S��9��!�!H�ɯ��~����v�7}��p�͙V�*3@�`���8CJW$���oN��m��r�{�*����ߓ���P��<�h�� ���N"o;΅h�{�9��477�
��O���H�N�A��oM��2�ID=���/L�������`@vٮ|g"z���ޚ�wDfw��;V^��8��< �q���@���X��ޞ�����󘗒c�~_D>0b ʕ��P�O"55��q�(=nj Ge�v1��t"�Y���TV~�y	����
��X����vv)0�H��.!�Y��[�J��ّ�o޸ͻ�m��W���226
��J
`L��H-?2�-��� �$�n�F���?6��{��ڜcֿ���ݫ"��k�Y��ח���c��">�o.a�74܆����G�*^���FI�: ���I� ���)�%*z����[�zb��yLv��q)�.��sr�ڣ����D�u]��\���� ��<J齜�U���V���hs[f}�S[[[�{f�J �"�,.Xs��tP\e��5R��^7���"bsy��%��.bN��"pd��hV�����;��d����\܀�v���d4A��\�J���߂�JC�#êƜ��j��o��CKpA��I�(�����a� �u�z�߮�R$���2�,���U��oP�%8��(�.�@n(?�_lS�B6r2d����J|@?X�g�y���!:E5I/�� c��U���^5fFĻY{e���'��?7Jۯ�r�
���+�PA$��B1G�t�Z��=/�S�m/���{����jO��%��M���9�v����7�V��N[�����f�I፲�ļ�dS�ɕ+��������G��bY�njnQa��i.�B78�����O���24���8 !VSB����Q&����?���^ݭ���������G�mNڼ9�<@q&$|A�J���mYK3.���TRo�A�{Kwi�4���˕��mETVH5pV7UE�v�ӥ�¤P���T��\�Uf��nl4E��'�,��B�e�wY��L^B�f�P��+�}�w����iR4��^^�輯��<�|�B��.X�a��`sI����D��Ŭ �$���5�q�N���0�)����ɒs�yO9lώ�S���h���Yy9Pk��~qq43�n�a9Dd��?L���.3C.���ޅ^E������/���b:�ҰD�&��������骷O{�(�w���r��9�N?�}��UܫI̲� �
$8�S���`�KēiNc#��gW�~l̲ѿ��H%����)����V�U3��?����7_��M�HT��7ֽ��h��W�:��~�|-���w+.:�N��O<5�%�<�j�'(p��`�/�����,�q2Z�8S�,$u������ �I��ԯ6 �#�#�EV7{����o(=ۀvI�u�O���q� Xs�~Ă����MDN3�Ej�Z7]	b����`�����$H:�.�m�?!qC�LU�[��H��MQ˿#�nZ����'ݎ��+���e������u��7�W
�"��W-,�L򐘄]SK��ۇ;��:Y`锛F노�k���v��n���	b���ݗ����S�6x�V����O$���ĸ���W/���7,_��yq����TF��TK���M5�����R!{�x������i�O&�𦬉��㛳��E����������?-���D�����q�m˺p	`�.I�ɑ����4���O�$��o~�y	��9r���N��`5^��Ϳ�#ֿBk������G<d�dj����$�;*�M������	o��^��sϼ��-č�m�ߌxn �� }�4��l����&E�ͥ塷k���E~)ѮTE��/��F�'�m���PT���l�m=��WC?T�Q�ڞ�C�h�m)p;|�`\t�T�����aH�# l�"�%cA�w��N��K��r�|[@����Y�C:��f�L����$y��6�^.o2��JUZx�S{�����C%TU'��&�+G!��VS&MPoZ��� 
�4�{���W�w���j�i%)�m�#�����ߜ��ͣ����>��i�K{B~ۆ G�� ���`'��*�&��'��z��ojྸ��K$=�d����V�5YY@��5 |�=4L6pPI��Iqߍ2^0̮�˨��F�],�k���	U2����WJ���`�ɂA9Ř��jr�P�y]'7��wHu��^R"5��8�ZJAW.�2#��ܣ��>]����RO�-r�|���פ^L��cCN,qj�A��7200 �ٵG岓i��Q�e���l�55�G��t8��&�T,D�?!�FF��6�;�&�#�� ���*�B� B= P0 �()R���H:ե�Y��oA�bV���Ѐ��/��h*�5y-"�qy���f�������*��w�+�=�a�v33�|�7�8�bU?��n� o	�~p�V�y�\d���/8����V��g��8�R2�
��W��*5�u"�e%yCs�!�-���F'\��{�W��=�Ž��o^�jr�.��`�uC<O�wc��:(���$��W���U��9�J�#��i�Zd\g$6�8f����R "�n}�p�.Pq�BR3�B"�Xl!d%�U�[�~O��_��Dk�Ϟ�*��s�X5�Z���8Gf����UBos)�Y}``���h�w�С'�b�E.a�L�d*ں�����_7��}��K����m�l/o�$�
��!���_��˯��R��>e�{��Y�nK9���P�n���n0��0�5!��7��撥�GX�h��t痜���ז@�rO� ��ᷚ"*'��[:2�!�u�y�))�!�(�=��Bj���s�.���k+q�k���� W��D�B9ڏ��O{�G��'����ɇ�6�?�����_d� �&���wE���,)�s9(X�PbU���dvR��˹�R7���w����0@7p[�ՕS1��:IW�e���L���_�P��迅��%O � �Y��P7I`0��7��C��'�.L��� ��Y�����ߠAю�u~�e�m��M$�]���V+�{L��1�o��M�/���������I��J ��з��wp��G�ӟN��i+�c)��C1�����?
��.���n)Sb36ұ EYL�^�7��u���?}:Ff���������ƌ�wEՙ�'�Bĵ�dv�Q����0���CAU���V:뭔-�L1}��su����7�����#��d�RX��a���^���u�A�~���n�Ŀ�`�6T�C`����#����`�r"23�M
?4!�=�O�p�dē"�e+�z��'kNZҕ������m�Ů�O�\� �i#�%��J��M�_����ad/�/������,*>�$���
�-n]@�klj����o���?�n���<���c�k^����}��������{�D�/��>���0�0�<��Ҵ��<�Y`z�+*�=9���nAA��p�7-+)<�>����ĸ"�L�K_5��Q.�@��vu���+5�g���o�e��i�#e���L ����V��|� �F��Q?.��4G/IH����J�%`&ޕ�����'�%��3)���t1/��4������ȇݿJ���T?��+܅�#��Z-A��3��q		H��G�,���!�\���ᦅGA��t|w��Ne6�E�#�S�z��lFvxz�rH!R,b�n�J�H�hf7]�i��d�zۡ�1")�֟��F��`R��X-��Q�W�^i�96��<�Y:1{B�p�`�_��@ 봵�?� 2����sӹ�R��F���y�/"Т'����s��HGQRNN0z�eZL��'�����P�����wzI%�Ԭ_C����)��g�|A�ս,�p�	�|>إ����>5��6�ih�i�ȍ�Nb���n��.痳�hnn�m٤�IMJMe�|����&�O������(ĸ���V�K��<}0�h_�sG�z��Y���;�|\\d�u��;@&,W<ȢY��m��#�����9O ����C�����(=��j!*7o*荎gڔ�e�1=D�����^��[�O��-]�M�s�&TKa�[�w�$����7cy��2�A�ڙ֯4����u���~'�`�����7D@=��Ө�t0� ����P���Sdg?�d�02�H:��

�r�����rvW� �ǜ��APxT ��N0�a�y���HQM�Yvdڷ�����.W��ICCܖ�fm*�RK5��4�H��漉0b\��P.�l�/�g�� _ so�~͵��2���h!(��X|��$f٧������һ�ZSSC �"�j��>k���E��Dz�5t�K�8���z�!9i��+W};��Y���L^�3.�K��X�*��z����dɞ�lK����2�s�W���ՠ� �ǅ�Ї��%��Y��B����aoQsy�P��c������E`����|X��S�fޅ�]SM:�n�QϾ�� Ϯ*a<��H-����������@����,�i��v1{��Z��&���������OB�%V
�:�������8�i�Y��e��`J_��|��[v���|�P;��ʧ�Y��O�.��jS��UVH��]�1<p$�g�QdA�7$n|xq����}T�o5�����"	�?57���'��k��Z�B��Zʵ��"UI��|)~�Cސ�2ˢ;�=��ב����*��r8�3�s�,Al��2��$xv��-�YK�6/)!| n;y;���`SF���!y�3蹞�����FQ�o�P�Z$%'?D��c���p�#�|�[�,�i8��,�Z��C��]x0{��؛���'����8��3�2�!*+�V�H�
�wu�.��!T��A���Ch:_�|������7�C�v�X4����)o�p�ᶃ���k�"#)M�HH�2���"�V	�1��!����q��:(x��z�|k�͟�S}	���&��"�z�1p���������B�
�q%�/&������}���t?�	�v9]�Q�|7���F6���@A5Nn�O�D�_^|���}�z����+��GG;|� r/ bYA}�t���d�������>�k���B��L�������/�k-_w{I�b���l=�nC
�i��h8�VVE_䗺��qj��U��'|�ȑD���ux��XB���) �]�%��Q'�h߃"�ׅ��F��H<y!�vI��j����M����A.y�g�ΛU�s�A�[j�"O��Q��b�Ή�2���i��°�u��KTBߗ����B�?����Oɸo�Ƚ�����*�]15&�I�za���p��@\U������#�WY)U9VC*�M�!=���W0UF�Dxu}]
���C�\ޭ7ZJ��[��xIÆ@l"A�*k�B�c��M|FRe=be�&��Jo��'��J^J1���9S>�* u��X�+$}����9���J&7;�}<�����Ѳ��//��#���V��m�=ڍ ���\�eQz�c [x��~kaCe)E���j�ܢR�jx1��9�Gn�o���n�!�p��?�B�W,���D�j��o4��8�]=�?_��p��,�̄�D�dxbL�}��� r�%r7rBFi���2�YP�4\��%++x�3�b�o�k�vus�H�#���B�x�1���	YY��eDR*܉���w���:�_hΰ�GL�K:72!������o��7�4E��]�/N~�8�� ��.�_�?��z�1E�)Ù�_��{dg����ri��[%LŽ$��P�a�afH@�����X�s��"7<-y"T�����J��a6⸡��۬u,�C�A������#���O�<!))k���a�4�-0�L��T^�F$���"I��t��n��C�C��1 ��>{���|+^�Hm���,�@��Һ�V��z��߆v8<��Saɢ ��̃3*g��Y��@"l�Fi����𸝧,nuSs��G�e�I���`�,�Q���A����!����[(A�ȕX��H��Wx�Ȋ'!Qkq����;Hf]�	2 D��n~n2K����+.Pg�XЉ����T !d;
\��7��[:耾���
�G���R�9b�Z��smz����|6/����Ka���R���Y �� XX8�J��� ��ꅈy�u���}���	%�6�
�x`�Ӱ���E-Û�Z�{����;(I|��yU�N��5���i.��h�r�|9p+�'v���ֵ]L%Ԟ��3�įh41c�h TIii�PO����h�$����7ϳI��WAꕺ0�&C���>R��F��R,�9U�:i�^߿�M���g?E絿���w��#��E4yoģD!\7]�T7�-�<�(�1�=0���ȍ-(.���'�4֣ffa����������>0G�'K<`�(G-P�(���E}"Y�������V\*������.e�r��T�y�H�Ql�Ic	��V��i�(WF޻���=��Z�����[�y��H���D<iY�$kѾl�c�j�ȯ@E��?����^s��W��_�R�>�Y�eW(�J���%���d�QO;���������Oi�s�Ο��ӱ���L}dS�a��WHGd)F���+��䑂R��ʫ�FD�� �*��K;��@�8��la���hl��KUB���O%P��V��͸)x!ǻ/��4�r�"�pƦ��V��g� ��sɹ��ȕiA�W���;����R���w�.��ޢ%��Vi�.� �b3<S��')�����=^w|?�Cb�(�x��qL���4��4YZ�A-vv� ���)d}K0"
��t��i+�ۃ'�gsgQ���=��4]��+m*De�AU�T�7��e�.��р\��ٹu�h���G�F27���]��g��O|k�v��a~�[`�۳7A'�����k̀���-o1��21hǔ��x2/�t:C	�iR�G� 4����hL��p�M%���Ӏ��� �2.fq��ݶf��E�Dq]V�Q���q���dhE��Wl�hW��u9T�"#f�/�$ͨC�I�˴�(�n\�ع�Np:�2��fͱ��k��b��6��D����gb�h4���L�{om����2���|~}�q�yn%��rJ���

�_q�U<�s�rh��ܙ�������]�����w�"2�2O�"�o$��(J���"w�8rQ�����^��<=� ��o��r�P�҉FF���\1T"�-/���Y\r$[�v�U��+�-��oi���͗��+�,n�}Ob����h��k�Rpe�8-=݀Z�q�"ДJpX��zKҖ�Lk�

	aK�
�]�����M��E���?�+!|��Q�������z:�>\C	a��|����F�1\�[� �ߌ��\q�F�f���`�����M�	B���ke�n���j�����QJ�ѩ������Q'��zd���C`��c_+M��k�O�]����9��l�'�h�����|�s�q�k,�RO}I5gW1�QP���ƥ��Ƥ�T,(�0K�"!ʗY���uu"{���dn�d.�/|@t,\��.���
��w�gv���"�:"am˯��Q�u얯��Ă��7-y�Ѯ��4�|:��k׊�^9T��M[��9�9�h��]���<����k�VE�.��V_k�w=���s��"m��C�i�i_�o��2S�IS����י���Ɵԡ�_��V�H��5��ٰ%��n�ꥯ�Z3Y��ьށ����\��(Ϸ����f*��[���n�3'hY�����QVsD�);�M��f�<����t�2i}�4�Gr��#+f*�gT�Qc&��*?

��Xrl�%Mg����ʽ�c�,�t.4����5���� k���M�]����ў-��+;�k���g����:�}���4$7�[)��P���:��{�T�`2T{a��O�1T�x�4N��fY̩��֦��ϼ��^%�E���������<k�cF0_��A2�C89�ɉ�y���-l�ظN��1.�olnv���k��U�&�Fh�Z��`R!g���Y���`��l뼷�Γ�Ƭ6<:u��b���sJ;��=6�p%�_L۴��=�Wzyv���0:���H#bܑ���&Vֹ��4d�>E�?c�/(��DB�x/��ʽ%7|1M��&O-�U8�ƲV�A��'���&��7���ivx�Ѕ�{ 3��[�Oen���1I��'K����HK+��QUn]�]�,$���?��7E�y`���7�,����J��~�t����������͍��ŗ2��1���y����u�FC1�:�{����'��c���~5�?l*�9��!�DpL�W/)�|�N����`��Gw-Q�f�T�o$�w��ѐ
�ӧ+-���Hs�!����0���E���󎮏#�feeᇉ�`����NN�-g�]�VW?����u	�������j��0s�Cn���V�	zY�,�ޒ������3t�#�_������,݄f}������~�s������c��/:Z���y�r(��������:{����T��|��k�!&f�Ċ������m��V�~�-���.��)�U�=>u�DՋ;w� �T�F�� ��
�sL��$�흛����������oު�;�󥵛��ieF)D�8ў�'B�`��T�8/����XzP	��8����6��h�2�58u��2�
=������ݼ�u��^N���i=��w���� !�#TN�k��:ȆD��,�����MT�"T�k݄p�Uf;�X��Py�YȐE�)���(���<M��R����'-�`2 0���`��J^2Z�N֒����鹭`��W���o���X-��
!%�!**b}j�f�J36O�ut���Y��T���7p���Z��\�7���;uu�<�ǘ�>�}�"��d4$�y����[H�Q���P��ezkh��h�1��u�\��M�e��2+�Q'`�rL%7��[l��'Y�=���wp� �n̞h^����G�u�Eut��F1*c�H1�(E�� �(J�"�� RX�^ņR54�Ra�.E�^E`i"�KY`)��ܻ��|���{����w�̝)�cd��W3=�f \����JR@��F��Vr{ �ˏޞȃ�F|�_m���qZ�V�SQ�:�`L6�37ڂ���w�%u��뭇���Y��.'�bHv�-at����U��nw�W|���nrQ6)!b����ݽ�y�J"�5��&;8}����Q��P��4��Z��1Gu��9< �9� �W�c���!�D�b,A�} �b����4���].-e��-LO��0�vZ#� �o#))��2�z>�]�\K
���r� /��Wc��m7�+q�"�wpvfL�y�U؏"x�zl3ei�ee���;F[�U�U�����|��i���R{�������NAy�#OMo�����5�R,N�xX��$�^�֫>kщ���Q�Ϋ4����@T>� �Vr	�{2匈j|I R��4�r@�EH�5p;�_��
($17�nw���9�-�Dj{�~c�_��ɖM0P�ج�f��)���nt�R��y:��]s@(dW�>ή��w�}i���.*��'�F\T�j/�z�Nl�,���ܐ�+� ��	I�{�\2
��&g���0u}lsn��T�e���js���>׶?�M��[�D��8p�;�����z͸o������&��� �* [�u��7�5���9-퍁�%�SQ�DH��'��)==�x&N���:18�ޓ���ڶ�ኇ�G(����ӊ�w���������U�M~<6�ڍcQo:' �n���a�0F�6�\�;^N)7i���a�M��!�:�5����/	L:4���~���X�<�_{�-h�;�h�z�`�l��ԥ�ը�����%,�W�?��Q�cSdH�}z ��=@A�[��ňX[����S�p&"Q7+�
p�����I��Q�Z�D���xZi_�z~��%��� w<(^^�i��Fx��J  8"�f $��,��'S�ǪD���j��d`���֯�	��b�Q���0�P��?� �J�H&�E�쎂��j�_&�Ey�F���"m�ѡ=/���2�y��\.�I�#60��̏c�G2���.yt����E,�� ��(d�j
8��#�p�D16���G����`����ޱ��GL�v�W���DTk�9����?Ⱥ����1P�S/����Ťo��2�5�Y?t��x��~�mX:/�U�=x�69Jb�\�$N%�
Ċ�(B�c�4S���C���G�����l���v*Tq��T	x�*V��{�J�	�0���L�f �=T��,__|� ����,���q#v��ΐ˟^¾�on�; =
��<^Ŷ��Ch�@M:<+��*䊠��[Qa�����%�*�'�;`܌�B�ؐ��6���]t��ki�;H�9�9���z,��a�@����^���z��~z�	_P^�t^d�F t!߸����3~t ��rS���['g�V>��hv*D��BPO})t�J�m��s�P%r�(�x� -�� ��N(ŏ��q��}2+�v��%B�BK�����@X��|��?��_�K��p�%(��=�
�D/3U�h(؀�Pmv�3 :��F.@��G�s�-t�ŵ��ʵ�/0�����y� .xTe'�},e"aw�	�������������6������.��vV���!�4�L[�L�a�!��&O�nG/6�<0:���g���f�}�<��z9yoZ�2nk��F�+a|w8~G6�c6)�G�u�<�"˲�0�QQP3W\�k\N��+l��9�r�؛JK�GOgI6�F$�!�E�(���w�ϖ�2��>�� ¾�R�7��!Z���xb���*��J���HN�C�m��=4�����E>���NA>�y�MXo������ �BP7^�>~����'pѝ�6�����]]	�:k�kH�P�J�zO`�=��q�zry�����6��!��S��Z��GN�����m���D�ku�L{S�$��S�v�`8g;�1��A�7�zR�Q퓟;�����O���Kn8!�d3��E��^���s*o��������`Q�`@��G���C������#W|
85��OZ��P|4�
�c���rP��S[ےl��h=M����z.�q[� RֺT��m�o;o��F�ah0_���A��oT�:w�X[F��3o��AD��7Xz%�7
��6$�=5�R�^d ׎E���9���+q~tC��$Du�E0��
��Զ�����Ц8ަ��oTP��|�M@�D�^��CN�����5��M�w]� 2�`�g��x��ax����(�)�$�����_� �م������{�aVݾ���&�9x�"P�	��S:��VOp8�̃����WIT��C�˲yqd�Q����\^7e�H�E��[ͬ@���ӥ���wN�3�;A�c6���mb*�۔TO�@ �������}^�fSU�LDe�cy����={G,�� ��c����I� �[r�1�n��9Iϰx����*�8�]��.�q]�	�|xR�c\��A�3��׬���2���V�N>�F?#���c�06��!��j�����c�ZA��{�G��!ѐ/Ҡc$���U��m,4
�����=�¿�h��34!�"��'��P�P���e���#������������q�$�W�2�.^�:��	ňXR������f���^�[*#�����	S�� &)2���/ρxF1��F�� ~�M7�Gg��n��x�mj���&"�sbGs�}����*���߶M�%,z7��5�)�W1�X�>]d�3�.���Q=%?�J�; ��p�"�[�\|Z�p��#�F�l'�+����xӥD�r�@��S!��A���]��czR��DJoQ���َGٸ=[����|ja�-�C��D��� ���W"�3�2:�5��c��3$ :=á�j�� �3��Մ�g��@���b(�LԶ�<=����ٸ�%�Bȓ��[�tZ��&�*���DoonN�}��b��!)���c�� �6���0|�����V,�O[G���X�}�Y�S�b��	���{7�6�Ю�8�cF����»�l,ԍ���t?`v�����G�'�A���Ui���e,��`*\E��<�@��/�;>j�PN,�4~H�SV����dC>}�]B �M��R�Wru�	x\�Z�Z�F�@��c%�E�UP~��F�a��:�����Uos� �P-? C��S~�C��l\�(�h�y�ײC |Oڱ���mA�n���x�>&����%�y@�Y��}	��A=݌����a��9n�����'�'�6�i�&2�����V����47�l���a5�̈́��D�;��#�����y�I]6Ρ��$�����F����x!��w���S���0�4������)�/�qd�N�FJ_� ހ���s�m���XL{� cZ�qy�+�/�"�VJ��}s����MT/���	��v�4
1�q5��t�8��vOJ��~��Y$*&5��A8��I����P�������)}��j|�[��ST�ȿ� ��D�@[hQ�� �c
(~Xh��&? �M�?�$C�!����&ئ-�혗(���V�r�j]��\๼��Z����Y�,�B�6�!T�Wb�~�8Gao�n2Aױ�ǧ$��ۭ����Ș�/���n�-cv8�s�h��J�����������Rj�l��C��/*���>�;ji�j�>����I��M (*n�+/��GV�����^���.��5v������^f_��A`x�G�%[��v��=�Ї�1|[bX10�.�ur�Z
rJ` �ʫX��K��������i�8�rA�: C'��D���*RT2�#��kk;�\��ޜ\-������U1�'8m�����ѨY3���}rH&�N@&Ƹd����`NW*>P�'��$
e�urU��mRz�t��:u��C*F��a<���s��m�:��#z	�^b :#���dol��h	����:8����~�J����a0��V9]�+��2y�4#�Ţ,��Y�$��[A���	�Z�����4a���kA�������B���33ڮ��/��"�h+Ȭ4��w��W��x�mwP�v�|�'��a��f����BxU��p+��NN	�d����Fp{X��)�����q4�bbx��~(�����P~,74�Ȓ�"�q-�r(�z�r�OS9��h]J����g�iOY}�O��Xբ��U'��ɳ����2�0����F�<%��1�����Y۬y	�#&s-�ຓ0Ћ��}6��t��9�1�������C�W�6n�"y냱Z�qۤg#H�  Ɯ����Yn���`�2+��� S��3�bj.��d�B���f�z��7al��>=���b��(��Pu��"M�o�	�μa��RTq��*o�vOG��妍���"��NM,�?��ۯ�EׯJ�6@����
`3a�`{#���ް�l�| ��ڳޛ�u!*�ʣ'�h�p��1ٲ��A8��]X9v�4.놧�j@�Y�΅�Fο���Wu����]	�6���X���VS�T(��ܧ�����Y�N���m�C�~L�߂�%�%Zo��H����H��L�dX�ķ8K���}7�n�C���\�k^�]�y�mр�>|�X��(&+�H�� �P~���|k6�׋����
�>�ᬄ�م.����>[�:]0�4n.d��k���F=���%�����	�X0�!N��8|-*��nY"�Lfe�/T��٦�!թ	�'�&g~!���}�J��8ݎg!�o� =���`J6涖�.�1�C��eC/�(gi�|�Ri����z�ꉻ��o����d�+|���o�	"6�L��(�̻����J[���^\��"��wo"�
O�R���˧x���``�i�bY�Џ��r�^x{��
H��[ȃH����	xC�k�e��v-�r@2��t�|�M�~�����i���q��on��t�oY�,��~�睅�8���H���L ��?Ru�@Ner����6��2V��#�&t�� ��j�B�O�С��"�)2�˧�5�e�B�ʳ(l��ͯdc���,�����;v���o�,��k/��6y��B��0}���~`9%��In?h"fU�@f&:�2���L�4�z�������h��&�%<�����\����*�!`T�Ȩ��	YD��#xL�B��yc��gv焴"��+h��zr�V���`����
�[u.���l��+�
?w�̷�̫Vb�
Jq
��MK����ծI������F�O�iH (�MH`���r3L�:wS:S~f �jC7^����A� {��q��PJ�f�����|ł���;�a��w�c��a�� ��J��R��[	��W�(�F���6��.{.��F����n>Xh�M˥�)�C�1�f�� rVrr �[B�AM[\XN���R� 1	��i�oy}7���Y��Nt;Gx�I�õ��m�����g�>�lh���� 6TI���ۍ�Ehu�7D0�����;��"v*����B"��)�5������	&��+,���{9q/I3�����އ�/��V`��6a��@r5_O˭��I}�{�n�^�@�_�<�Zxj�R��N�������(���}�]�<6Qu}�~�����c�D=�Ѐ�8{]�l،�/"���X��z�P2����h	Ovv0	�q;L�ݥ;W�F)9s������]?�{���&��^+�2.'+����¢ʁ��-oz�})Q�WJ����׬��/�F��2e�4&V�FO�f��'M7%\0�d��ؔ�ed�6�誂�cOS�a<���]9�XJ�T�x^*/ ��d/�
����t�b��ls���6�g6i�;��"�y'��Յ�=^�$�fp����v����ۧ�`�L)��hbd@���ꮔ�E�5�e�j/q.�V��Pd@���a��8�mr%UTWl��$�D��������F�]X�x
�R&$��z�X�����$Dૼ@ �~6x(߹���c�(���f5ɻQVm��!�(T���"zc]o,��������&R��b�zϲ�U��D��Y��Z��К~�ng�FS�S�����+���(���&��F��8�%:��q�K�.ho�V�������\	�O:�����6�x��Z"�+((�KӀ�J��h��Ou��>�<r�"j��=khcʣK��S.(�FG��������+��n�۰�8��zԵ	�]�y�����Znn��j��-�[.�jw�F�eN}(������WυwD;,��g͉�+s��5�H[�#���WB����!1�{��/#:�L�9��c���i���fz���n%s��o$�������m��=��.%腣n�S���-�ߕ���>���@/l��]�j�<l����;x?%V���$m�z��]m�)խ6yPtD�S{���{��&�9�1M����t�G`�,Y�1%��؋/S�Y(jJx��[|.I��_c*��w#C�� ��b\jʶm�[��`I�N�������N3�����h��Ѱ>�);9}�2xכ�[�n��L���T��������m�pJ�Q��4>t�����iW�u���Zp����e�O�>o	��;����>�*�I�'c��tf�{�>��H�����n�|��w��������/^����^Y�.�	[+q���41uV���(c6ЯVJ>�u�\��8\6m�Y}#���۲�F��%�֭�����"��5�[5� 81.~0��t*]}��낞K�J�dk���$*�8�;<{8H��KDҗ&�i�N�n�q��Q;n����q���gQ�aF>����i��$�<��ކ��l�./��N�;]��~e�:��Ʊy�����𳌇	^�y�_��4�I5V���u����8�=�T�mQ�U=gN=CY�\F��&H+&Z�%[��YSq�zd���/t�����ꗹ�0�O�����k�~�.�;oE�٣,`�p�C����}ʞ�!��4/Mt�4!�[j�&j����CC�?G�
~���Qd�e�z�))�<",.���C�1�-@=���#�����Y��*�"�H�c ��ܶm(ى��0@��"�T؅6�0¬����:$�y��q��>��,ا-q��ˮH��f����z8qdC;]ch����!i�Q��@�qg�YCBB���f�̧�A��#�s��u{��@8m��z�#�&(p7�|�t�]����� K���=��H+hÌ�!M��2,�x����g����I���2ܶw�OP??���>��U'�c��f��Ð ~b^��Ky6
?�P�y���)�{�,�UkƤ� e� ��5��.�|��+zj�MY�hw��|������,�z��Q�!����s4������W��.(�]���KS�˟�7�v_�f��o2�f�T����%ϻ�Axo-�$��.Ι�n�-s�"�/M�e;L��ͦ���+A��L�ժBDAT{U���`
RK�:�����P{^E���7ڥ��(}Y>`դ��^�'W����Z�e�`��r�������ǵ��A��6�&��`������H��!J檞S�z�&vL��^9�&w��J��؛���)�FOO�,����ƥ%+�eJ�����g��Oc�q��;|C���|�2N��o,e-��3<�܆�����#���:�����r��J����B����T0���O�u|�
a�\�|vM]����x��˶�]1�'V�%(��Y*A��ʕ���n�%b���v�^}�9�ZY�Z�����?�#;�W2�G�@#5`�`�4'�/[a�O�Թs�w�Ǐq��W�h��#���$7��7�j��	�} 5���VO6��N9�`�m���N���32����vl���˗|Td.;w�����^��<읱�r��:���OXT-V���--߾]u�}�8�}?E���
�y痧��~��-�?,�D��C�`�=x35R-� ɇ�ŚJ�Bl1/%녇��x��ִ�����U�/����o�y���"'��^8���?�����f4��<7�~8v�3L8��r��.S�~[QJi�{��K�ю~θ���s��0��~�0h��B*J�*2�p������.Qڇ�o�a��z�:!**2�o�����Ń�ū�2/���.�߂?�=�2U�2qc����n����DU��-��ƤܥpR��*�n^1A����Oo�j9���W�^{m�n`iްM������s
K����G7��*�4ͽ9���K" Tg�|	ʑ�6YY�˱�[�;���h���Q�9�k<@����d�u��҄5n%���ƻ(��mch���h�p`�9�����Q9�LA[q�e(���O�epO2A��0!n�f��8~p����[��P� � �A��)(�>��o������=N2��"�/���Ԥ�ƅu��M�́O%Gy�ρ�5__��<Vd�溷��>\ER׷)�J3ٝ�Ln�m� /+�/N��#��A�qV�R�%$߇]$GJ�7Cl���<���h��<��B��
��{��u½|�g�j������u�w��X�1��_�F!x}��[�z�����K̞�: �y�" �A��ƚ��@v�JV�w��+',� Y �yfD�!@@����-/���l�
v�F��<���VnJ�r�({��B���C3���Q��o#A���J���������X��엡ܦ̓�䚹9�Pu��i��˗A�tt�ݗ��C��1�:J=[���ш��Q"���:���N��E�$��6�j�xe�����2��Q��>J��	��/���7͇�q����@i����O"+����oHQA�#�����7��/��U.1(YJp(V�l��]��G��!b���3Z��W�a�:��	�C��.
����_��������guu5$�P�֥����qL0f7��8ߵZ)(���O�̳���P+���vx��ƕm�x�L%M����fR��&��D�xȡ\y>���KzO). �Y�z���N�z��ϟ@Q+3�A�B��\t4�V��n�r��'f#���]~B�~DP�A�8����!�K;E. �h�u��&�Ck�����[%7�j�ع?c�Ƙ���zf�3�x>A�g�V-Ŕ s �o���\/�)�p����?��Ck�z���=��̒���ȓ=��OIC���f\�7?ko׋-�U̏e�|o��U�tm欤, dv��;�D��c:hL����	L�;�B֓�C��1�L���%m~�ing'ũv�!�˿���@v|�e���Ok�u!��9z��xez��h�JxD0�Mz�.�u�wƱ�ޡ¼۴V�,���p{N3�􃠒ݻ\{{8{�r�Նz��eo��8�;��e�Z����[�2o_���Lq�\m���"��U-4�I�ݞ`j�S�8����m�����is�֜��g=n����S���7y����m�G�2��&���ՙ"�K��)���?�n@�W���ya�7��B+ֻ�KWG'{��� .���DA_���[����O4�< $���2O��#���-Ŵ���J�k#zR\S�r������O�78�Q�)��	� i6�(�2�`J<���Vn\���=2�8��7Q�#cc�a��"1����{Z��,�Î%�H-��T�j�#������|VN�s�����=�w��ۅ��֌�LԽB_8��NvL��<��+��;�!�;'��]Lj��}�,� ���a��R�R0Hy�}��maX+7�r�[h+�,rw���Q��{��nY�.0ԁ��|LNQ+�N�c�׬�.��i{{;�EPq�A���W��CqO��������{t�8��˱��kv!��P�hZ{�g0�kB�*�&oNu�y��� _�.�Ր7���SX�����Լd���_��r�HuR+돷d��	>�2�ڡ����57Q��$�<F�@&7o!4C&SM�Ug�����f�.�Ⳍ�P�ڊF����7��CFq���9���e���9qD}Kx{i���[�{�\�C��"����~W$�Kʷ򅷓!���\���*6['#��}���;lZ�ӨSJP��N����X�y^�&+�QɈ�f��@�^\�"*�7�q<����wl�B^����Ug\�: {�ŀ�{(8�L-bv�:�"*'�����LE=����2'Yށ<U*�:8سs&�	���/��S�0u��鑎�N�4��;��+˯�q<8���R�T�mڀ����R��e�J�C�>5�D/��;���:e����hy��0{�:գ��Pٻ���]� ���p��5wsC���]cR`'��`_�l�����;����;�ĝ������L:Ȇ��G{e��j�_���9�d�^TP4�<��r�I��aC.:���u�6�l�g�W�K*t�RT���v#M��1c�h)�<�p�d��k����0��R����'�,&�!Vc��F��a�\��&�Sa4Lk�]6⎅]��|�47I��:��i��UPל�y�w����];d���4��L�8���Cc����D�Au�ڧv��/R�&�X�J붞�l�L�t�P����%XB�l���(������+)�uJ��D5�bf���SB��K7�ߺ�n�7������ݿ;�Y裭�JroW�Ā�Aŉ�&������KWg�ȆU7��'�*n!��:<ِ��yG�㬴��N����7���S8r"g��*��M-LtB����WPJb���OZ[�����Fљ �ߵ ���|���w�R�}<�~t�
�8C���4�=q�h�pP-5u6 ���[��ؼ�E�[�PPV'�bH0�Q��R�=mȱ���3P��D1-p��� �ݟ�r�WW�����%K�v+�X�z�:10�6<� ����$J�*��8�ʆc&�ݔ�#��1hX
���"�Tr0�y�a�6��f��r&a��� f|��`c��VE�X!�۴n9�95eo��_����$� HCb�?�sB��Q�.N<��;%�dw���d9���o�1�nNY-�i�w轢�o�A�OE��=����F��k]�r��<����� ��N��q�.=�u��l��YB�ؗuho;�~eks�*�F�J��2q4 U�5'G�&���N���b%�3{Z�~�r������4~DE�-yX��������- {dd��hz{�D!0�w�l��L�q���~'_�_YA�Ǿy����'�U��Ӛ�/:&6�vȏX礆�'�.�'KWMPL�g� ��'�J�F���e}����㊡�څ~������3 ���x�n��Zr��Lo��OY�@��Xz̷6��4�$�] �&��
@��+��&��Ç��e�l����7��gfϞp+��Rl�dl.��R�I�wZ|��������31(�ʋ�;���5�"_�D.i��w���#
� ����f�����]�I��_P��:��xnC�o��?�Ր��rAy�"�W���ݧw���W��|��!" ��%"֕*�m��L���W�7b� �)��ĺ����.���- a�蜑j��n�zDn&_,E�3_��l�v�tu�Z�,*|��s���@�5k�C5�]/A��(�U:~QT5��9�)����㰌|Z�60Z�%JȠqWN|��T@�? Z�;�8{��K�577����UjQK��U���/J����t@I�UN��V�%qz���)�� ��(8Y���F��..y���<� �ğWe�׃<.�(�M�%' Dv+$�p&j�����r�5�MZ|"�(:dȝ~�e�/rl#��H	�����0�+�f���&���.��CՊ�5�Vko�Cc�+3�Hy)�{��P}]��h�R�b�j��.���/\#��I�>��j�bd������#��@^',K������㦓qg�l���_�Fڃ�O�F� �����luT��O4X(�es���b�Rz�K꺛;lӨ�E�"���|ʸ��(�#V|����[=v���Z�-��۴Jx����E~K���e8�\�{;�g]��c���Xeݠ:i��_�	7Y���D��:�H"�d5${v����[=��xų�m�kЛ��s�m�1_dL�*����f9 ���\�(ˍ<J~f��띜W�ٿ�*�oF���oP����4ǧbګ�����鍊WL�ԸB%��p3�_x8�����q����x�fF��{�8���ݘL�=�Zy6�VRd\��!2�i߫�\7V�ekM�|ƣ!�2�b�^��T��[�tUu�� �TF3��<��{۽�r�]W�?)=Ǿ�wdⳡC��W�k�p��ʃY��e:$�6���[]1��?P�������i��.��X:�} �
�^}tN�O�7��O>fg�'���؂52���4+�b�!S�x��z�/� m�=Կ�d�)�;�' ������$��^�q=�^?�!A֞ȒL�l�ך�ܷv�%ߜ�;�x�/UM��e���̃x(��(w�)�' �6��� M��&��Qm��Ǘ�[��U��Y��Lʞ����'**���v��k`n Z$����T�ou�G������>��g���#ܭ:)r�V)�vS�G���Hާ��)���+�,S3ԫ9�m���^�쾱� �<��wCnl�͏�K:�����BO��y�#r���@ x�G4cҿ��KoU�M�(���@�x����`rt}�ۭٹ��L���c�0��N��R��k�P2�\@$>�hv�4w]�B$�������!��ׄ���&��m &�6Qsj�0N8���<�89M�'L�i�g��1/<x8L��B�/�� �QP�:T��@֫!�q����W�Ѧ��n���5nP��շ�T�e�K���� P��-��3|d�/n�1C�<b���p5B�ox�?��.#�:�7'�O[P�{�K�!�F�s����d�0X�4�4n�F�����S�Es��d�Yy� m A�����m #��x2죈:��YkE�l��Y򶟣r�c4�N�j�ơ�0܍(U�b�@�:be=�8 km7~��a����z?ȧp���	L�qBF����k�(� G�fK-��Afhj_�'Yq�LoP �=c� 2����&KS��2�*�{��������M�	0��T��0��Ғ�� �\�46�פ�a�8���|R�a��mb��2Rjr6S
��o�)�_��Ю�TtH�������-�mp=�ybH�\ ��7�+UAa�`@���n���	�i�w�F�Ͱ�O8�����[��h葻���E�^_$�����ט��^: �rJ�Y�SG����rN|��R�C����w� �j3[4i�IU��ܞB�GDh��E["��V�|�_Je�A�Xt�%�͚u���9
�|_��`�Q��&j���-�NfI����'����^��$��@��w=�K֍��S��_�,��3�6���u|��a{�'�}�u��ѻ�e�̉<b�1C(b��s�m6>2[�Vil�_M��9��	<\*Cy��gUP�d��@�Z��^|yni:��j7'�i`��|R̷ɋ�\�@	$��Ʀ���X�o�K
�Lej����OS��1��y�X�E#,>��y���Zh��O[[[�|t�ʖ�zĩ�o�;��7���ʔ��zES�?j���#���z��}��\F�]��L��FY*/�G����� ڂj�$==���SP:G�G�������ny��7R�K����M��W��V� ����N����C:yS�<wG$_�Z)Tn������"������Mn5Q̗F���wl�"5�����(�^kd�����70B��qZ�ܲ�a�T4�)���2:��rj$�KB��>��/
ܡ��4u��F՛����/o���go�O�9 �T>��A����i��U�8Sp��0��iW�;��_��y��~8|�A5�l��8	��'�)���s��Nj�ڍ���|�SF�s�Mޥ��'���<n0[��N­����!�uZ����1���(�e��c��+�(|R����J[�������yൈ�J/�8;��ZZ���m��p�68hG��3u��@��0�	�E2$[�I&�׉�g�q�4(3j;���Y@ПVW��=�
�h`&�B��
����D��l?�]X���G��{��
��T�*Z�=�d����WN����e�t������rQ�|~r"1�Loy4��Dz�4�Ɵ�{��_I~T9�/:�疝0+Ss��`g�Ǐ�q�݂�a�@�U�@��?�JCí�x���1��r\Z�za�Z(��E�����L����%�̠�Fض-9Cv��փ�_)�oLZY6t�2\yd��1T��F���XH$�.��k}�c����[ԮK}<���ԤYuS�;��-�9�
�#��m��j�;p�۴�R�&q!m�Q���<
S[��*N�ӊAx�Li~�-�*�{��O^��~�\�Fa��O�&��� �a� ;t�CU7��5w��91{t�fB\B�K۔5/��1)p�����w{�6�����Jg`��^iud���Fݶ��R��3}hJ�%AOl@�介�S�ܜ�����Ef��7�L����J�B�P.e��Õ^ �;P���B�CIm���se��Z72��!������"�'Y�6�[`��rs}m��V�n`/���"v���]�U��Y��xm��(�h\4}::S�>j����9�Id��(���i(Ń`:00 ��
�W�/�_����'��{S���y�Ά��{̔�����qބ�����`�r��>D�q���e%29h��^�a�:�q3j����ԯ�V�xv����+�����P��e~(���:�b��˦ nɆn���������b��뺷�ˤ�$�j}}s��DS�
�+�f�}��q��p���c#��\r^��viD����S�����&��A��T4;�Cm���A}�x�����߰딨�F6Lb1_���y�}DͶ-�GK�¶I K���v�"0�@�G�PBSE���T.�	n��.mRt-$G �j䩟U�ޑs��������7�9ܭx�<Z��m��A�^Sw�_,s��'�-��F�i��@e�m[�Fx䱟�L�g�s��s�<���r� ���B�q?���w���M�6��#��/h����� �`G�N��=54y��������M��Aզ���g|�z�c����%Wd�I��3�h` P=ؔ!n����_��)TZ���P@���v���,Lt\�<.��w�����f�
+׹aq�|���z����[:b�3��R����F�9��)���Q��őZ�A�;� �(,8g�~Ě�CKV�I�yN�p�����^Ya�Ǩ}Fjx{{��f%j�����H��z���A2��&pK��D�+í̋��]���¦&r�k�P9hR" �j�T"W�����֞%鑐�?Ev�.e��s�5�ޅ�ل��-7
c5U0�6�m�ݺvݚU���{u���������9SC�g�	��r�(X������Xxb�t�;A��+�b%�f.���N��q�g��T��<�*��&**)e�<��+P<'��x4�f�N)�������3���@�I=}���m�f�۟_�ȟ��CG�����7�d�uW���-����",�S��G���9��/i l<�GTDD��62���y}�wѶl�!�.kKC��7����
��_���N�Ww[��+z��q��#���'�J���� �Qj)���C�޲RW,B�׎G������^\~�*>Y�*�zo>��u
��-������K�0dＯ��+��W��M7��.�_D?+��z#^FG@�r��r�����9z��nSS�v�S�bRW����g!Pb��L+�).u�6��K�=x�D�7��4n��P�k��=E�����jF�#�ժ��$�=��ސ��#�d��oViT%�]`�xC�RzkU�Ű�l�M�tN)QF"��٢�?�b��e��놮����?�rA�/0���hd�?}d�A ����s�U�$h߆$s�im���sB�c�⩆�S��J<����AHs��kR�㭳���֖'��Go�u�ͻ�C7�|7�<��u��FQQ1AG���	���KU�(8fl������B��*U�![���)[D�����~�f���E�MU�����l/��L�^�G��y��%t�]<����)_���,��0�޵�F�;�Qq�En��::YP\�mc�<y033�lRg�I��Of�`�pO��³_�X��@�����M)�8PI��U��NB��9��Ř8%C��v�yaX�6�f`@���Sn�/��NjpO8�X���X����}a]�=/ܐ����m�����ݫF�ۼR".y|�����o�2(
�Ğ������@�ߛ�1;��^#�D)���%[�EV�漩�K@?�G�vk�dK����{�5�;?��j#�a}�Ő������C1�t)#rssӥd~HI����.��y�:�>�_g���%f���.�v������~#��A�~�-#��pC���x�\�2��� ��yK,�<��*0�W��B�D�w��K*�;�ϻG�>�r-���<	�AQ˙[֯:o��;Ք��W�1��5wAc�5 ���k��kwq��rny&)�4�#�xS�0�)��k"�;�nu�$�
���e�����ζ����g�l�4
\ťL{�M��9������E�/�*���b�cR����[1v�Z����*�|�w�ؘ���>K�����u}_&�*��w�jxxx�ٮ;�/?ž?(ix�n�`w~H��_�����Jd��C7>h|�Q�jr�4G�Aː������Ðf< �|��x�����q�#$�<���b-�@��U{���&�g��'�Q����X������D��;'���4��K
F���R[M��hgx�s��u1�F��,��7�X/z�]�
d˧jP4
Xg�.��𐮨�D��"oι��V/={�Iq lޏ��:���&���/�0}�_ж��� �e�+��-��6\����X$:�s�-z��#����&��L���hV��fo���>R�h�%��Ee[�0�����D��*L�۹�q��:gay\Ո��n&3��S1d��b|彾6~�J`,x�ȅ}]6_v����ʴ������5u_�
.6@ GWI�A*Z���9@Y`�Df���s��1��ͯ���v*l�#�໘H��]jU�;B�V�Ɓ��UMyo�,r��Ï����@6nb��㮱k�Nj
�S�S!>&nY�����{_Pt)�mS�3��o-.��7-�E��k��q�Prr2������u@��$�Ҍ+_��M/���@6��\鳐̇���z�އ�W>�`�Z��7�?�4���YΦ�Z÷�.]�"]3�5�����]�6�6x ��PUx U�W֝�O�<�X��2��f���2.oXS��Q)O~ ���FKk�gec�D���v��9����C�1�c�`�{�ۦ/�D|��+��*kf�B�(� ؒx�<��̘�:��*�W�#?R2	�tx��zɯ�˄�=oo��Ĩ�����4tIv���1ј�C,��X��~{�\�s����1�@���v�����ݟ`^t4Ee��G~�n���ZU��۪f����rt�3)�q�e3@w0@ � �ן����FE]�T6��͜��� �]aQY�Rr��I��7RŻ]x�k�eA�q�<F�zP���!A҇��t�;�t��r�����:�i���l�u?�!��b����ɋ��� r��ҏ�=�0ԗ�O�WuR�^&zE/87��>,�&+��c>~W>"�5@X����=,��~�ر��W�~	620!�.@�M7�O�X�胸ۊ���E�^�WOpe��<	>'>u�<T5�5me�'%�K:<��2�����H�&dÕ�<�/Ͻwp:ɧ���~�B� t�BQ�U)��~�RO������1!##�����x�m���&�$�yP�ytE��W�#�}$��~�Э}O` b�B��h�5�ҩ�`����*����G����O���o�T�AH�DM��¯�� GӅ�;��i�����_��4�L�@��?����{���0�����H陪LJ������m^$m����(�(�������Ϡ�_	
v��ߏ�||4�2�i7�#�*�T���#eZ�ݗBg[4+��~E�u���?�;M��`��m5v�Qɟc�6`u��m�ԉNt���:į��t��]e+z�)t�i� *�1�3 �s1s�j��09�&�B����0XP@Q)��=��N��%u���w�g� 	j���w�n'�;�X%�ߎU#��������K���f��mn��t��ټs��v��J%�I� �y�$\���[�uc�b,��5[��4�2���t�/���~�Qq�f�y��ɖsF20BFa�'j�
J���iMew�%��6�w�զ�\K�1=��/[�Z�K9d=$�Sq�k� �bc��. �D��.�l�މ콹���˻ޭ	R�5�������{�3�:LR8yO%R�Vz��r����g	�	�#Wa�rk�^�ZH�W;Rs�`�~b�`n��	�[۵�
2��uF;�X��V��;���E�Ʊ�nǑ��|7����Kn4�0qx�2�
3�һl*H��8p"��#T�L��\[G�Є2��^�3Sz�hhz4}�s��8�!��!��=ExNЪi�dG�K�r=����1 7Nv����H@��uu��� ڍT�!&���ݏ/�za�T�q����u�&���9���x��CR���r ��ҥn��][С�|0��b�&�n�Owv��Kъ<i�
��C�lV4�_��nY��u�p~�10��v�L�P�Щ���q��n!�?D�@8��1�R�N���Ӱ�����P�@޷�����M9��]T2t���]Q�o��'z��,e��$x�6"���ͼ����K�{R���^��c 5�6��W����A�������M]�j�[�-7�W7N��F�j�Dj�{^�J��s��f�䬭KV��6��\v�ҥ.2D�	�Ni;>m#�L?I�9��nyOCHtPKu7)_��J_��9qFS�fF� DPċo[���v�)��9�N*�ZTWQQ����c��t�%�,��?�K*��v�%>�]-�E��{�s�L�l���w�0{۞���k��u�w)�˜�Ka�/37�8n�����_Ż  �{������^ߊG��եP��Y��Y�}nV�	��˽{�{���5��3��/�S\y1�����b�N�0E�2%���ۏ` y#��PT곑���HIA�4ȗu_�${�yy/� t�m�ked��I������jr�o:�JYY�'N�9Ȇ`�/B�>#��ư��p%|�x��Q��qYf[��p�����R*�*H�c�"!! ���� ݠ�`Q�H����t)!"% �t>R�����~���}��Z׺�����w{��ğb�/!3(�4L�J�rq@��Ò�,��YN�/��8��~P��+*��R�S���>������#���C;��ɂ+Fp��YN�b�@�U����.�]��0���f�$d��C��i||y��Z��`+ *�W �og`\u���}=_F������y3u����^����f�v��ϼ�V��Q�ٹ_=d#r��|d�BO/	��Z����$�' ��}�\���mJ\�A���&5U���9A��D���)*)]?�3ښ����tt�Ed	g �	�<
�B�ɦ釩�zƿ��6e`�Zp�á4���.�i|o���r�#]tf���uDx�F��8�\d���,L�P�Y�eA�ys�~��Ă�!^<�����է��n2n%���g��y��(��q�������k#���F!�i���a
����I~���*�U�.R>^��D?)� d��o�GK��aѹ�?+��dd���}���١i־Z�il�X��q�Nq\��'�"�j�����d�Za����I!�N���!���|����cB4VWm����Y;ͅh#�Ј+!��y��`~�Ҝ;u��C�օ�n2v��`�c �I	G��*[���c�?>]������~w�r쏍�8?�9P|��l_7�caL���.e��o1��hEj'0�$%���?N�/Q�W�A���2�
�
�:ζ��^�&(s�MʾfǬ�Q��]k�lԳ$vxK��9=SZ���Ņvj�q�#A �����db?����l�%��^U���&f%��+��x�a)��+n�cw����jq��f�9���ȱ8aINi� �:���=�������Ǐ�4�2vX��>���m�(���R����F�T��|pآ�c��<�\�3�5�<�M<��yR�M��|n���~_�����ʺ��%y@�ǫt�`e�T��k-���( GL
JB�&�ivL~�	:�k�vK�k.�^^�13�t�-e����Vd�^�.B�����4`"<�]��)���!(x��) ,5y*NB�9R���!��e͉�[L]��|��y�ӑ���滪$Wڠ�x�%��{��Hy��?-��V����u�Gz���_L����WڟO,NV�ʘ�౐J�sC�>x�ZPJ�hct9��fmm��f�� =�Ԡi�]�o-"�r��R����ț�'=�����VS��(i�H�E��[:L�����_��@�;L�c"�t2@��Б�����_�_`U�wv����ؔ��J�����<W%(h�U��]�����H̛_Y���$ux�ή�������/mY�ب��p�f������>=>HpJ�q(6��H�(�Xk7�V5f��l�P�Ԋ9`!�CBC�(i���̆��+O��f�h-��v1���]�9`ЛfW��L�#�\S�Y��]r��!��fO��d�;��|b�u�l�UEGGwg��WTq�A���hg9福���6��=_r��5<
�&>�9l����S.��g��D$�T�E.t�t����p\!���hcŢ,xO�R�b����܉@���Ts3��7Р
��V�M�#���Ę٘f��&K��^�4�k��۷��3Z�;"��즳�gk����m���ϕ��8�ɢ�4�b�����0��?��qX���uKk�9��!�Q1C\&J�`� �ņ9�ք����ރ���{� @��p�Q>�F��GHw�Y+
,������/4QSX�k?arD҈[��qa�='��G/��5����HT�O���y�\�\��p�` RJSEq"��Ȥ<j$5�|��"�{��o���wwR4�N�P(/���prFdoYr��$g�y����α��a1�`�G����j-D�)r�[���sK�T�����LWs����z��4@+��mK/���Z��k[���F��@S���H[��dd��������s�/��ݝ����,>ZX|=���̯�2O%H�CNW��*(�AHb���0�����F�Q:��2B
0%e%O��q����I�݊aFFF���+�ǣh� ��ўc�封E�����i+ݨ�ݱx¶��yp0���篸�j#�Q�Q{s�rᜆ	M/�'�.:^}�l���ʶ,�cslsBn�(�:�-�2U�L��K�ؒ2?��������8�m p�������.�꩝�����M����\�4�;6	kn99�!y�M"��S�\W��*�@@�9�o�///���{��D�`��DV��� �
��~�r,j�Z>>��m#ZePvD���,)��/����3t���0�E]$��;A)f;��K���fJRCva*�I�����|@̑����w9@l�v�{�,�^�=�88�K�en�ΰ|F���'�@�"ɲ��%�Q��7?�����Nေ�ѻ`��og|�N^bۯ~5���He��>lt��oNnk��V�m�=�\����R��@�'W�����UHт�r�|����}��]��옃K?�޿	���H���L��?�;EH5ygD�j���f`^��r�����I� ��uʯ��؏瑴r��,*e��I�l�a�6�nл�+v��46+&]��1@>q��Jڍ��v ;H.����Oԓ�6��I���~u�F��h���4o��+��il5M�f�u�"K
@4�xWS�a?&G!�X����m5�ZZ�������U���)���[x��m?׀ڍr��Ò���7У��|eh��TD��u�۩�g���L ���)�ݛ��o�iʥ,Q/'Qk�ٽ�E�CfN�N��-!YV�J��9F �t��/�$��ʲ��eJ�~xz�S5,��y��C��yh��ڰ$�dG�������0���j�\�IB�ל��tD{�k��H��UR2�Wh���-B���ùB�9��"6�;�d-s�,Yrs>�"-О��!}?��3�+�/�!H8�f>r.���w�̷��p|� ��v�X�������L�"_���B��;�v$������{�<�2ov�O[�"�����f&��{?�Dه����q��2�ha�4�ITc��N�k�]EoL�/P�A�bd�n�r�q�F��	��#�����l���/\����Of��l�)�� d��ȯ��A%�-y55��u��u�u�;��S�1V:�yO�9)��EeFd>\��Fz�,�b�x%_��<���wfH����|�h��3��0&ܑ7��H��l��`_?/ʷy�Y��Jx���2/cs����,I��9�E*�J�I�E_����� 
ncc���KI���������y`L��^��IW�L���}/by*F��4�l��g��S%����<�g���CJ3O�[Z��5��$h��:LV�Ի�W���|�tX2Һe�늡Cs����c��-yw%��,26E�:�0Ҝ�
��7��;*�	�wOyG=�!� k��OxY�-N�^ݦfP:?|���c[�QՔ�w�i������1B߂`ZmWD�C
#-=���ѯ�֓f�#�4j�Ә�~��&0�2$jd���"<�ԑ�d��I�^t�Z?�\G����q'3�e�*�uk��u��*E;=�N�6��t�����d�JnC
^��Lz�+7ė�����I��<=-e[��CǸ� �R���^ W!�V	feOpc����v̚ۂh\,��%�ڄPOz[��d�yaF�X�����	�zVSy&���ҝ#��gee6o+�-i����`_��ƽ�b���wwfC��������������o$m���X�Հ��ҥ,�Tn��')��I���Tr���&���ÝƲ��cR����hhtk�{���(����~ץ����C�ny{R=[=^=�\8�T	�����n�L]Ĳ0V��ba�Q���2�_ř˟���Ӛ�F�c$�Z�mLm??���DL����of=]E�a�U��09]��0F�Exz��n��ݘ��]�Fܳ�X��[9]�Wְ�����4��pC �YDh>�]_�XN��q3']7�`�옷�d�U���za�����con��Gޡ,p+�b%)���{�|����(5��ח�4S��G���c:?�p3��=���@��I1�y��f�j�?�8�$w7l���}+��}��G"�`M{]�E�cܛ4�
:�L3��L�P�A�q`b)�>.޷�a��Vk:S��\B�(Uܡ�E�DT���م�A����xn���Y�iۮY!���T~�>������	X�x��\͞�*��b{�!�z��!D��u�<} P����Z�;�-�*o#��#\���/k����ܘ�Z�!�X�*�GqY/aʑ'X-�x�.)'���?����Zy��,Xj-�f�L&u�ؑ	,J�F���	ׅ��c���
@4="u����p��x�ߎh���Ǉe��r7�s���ܫ��&��$a���1f����.Ї�UZ����{�ßo!��q[�u�Ѯ<���s���u��=s��
���NW-Q�݃F6�A��r�FF�6<ɪ.���߷۳�����i��VZޝ�p���M�Mm �/��Z%���?AA��}#�Wԛ���H�Y)`d�v�+��ӽ�N`/�p6h���ٔY.����u�b�r����KY�A���Ʋ�P�����.�m!�+}�$�h7��ܨ���9XៀqX}��kcN +�'���z�d��1X!��k���m�<��:PWoc��4�g���N�y����̡��9�k�$]�7���#Uv����m�j\W�^��,�JE`��Q�T�oW��A,���'�|=��'��ChRK�denњ���8� �]`a=�1��:������̗����������k߃�ۏe��a*�'���U�^��9�g?��Q�>aR�b�XYYy�[e;]f�M�w�ߑ~B��r�@��h�����Dc�������0��ɫG�_^&��Pv��ݻ"B��R|�B�F:�o�+q��e��O�\j:g�^��<[^�����/����'C�O���l�/v��Xs���%/�'%v�©� �啾�n��@y⑕ҷ;Nod$�ؒ[��{��Z"�
�X���3M��2>YG1�����#,+aR�ķ��]�P]�˅�����b�]E<Kwv��`�U}�폖�����]�ew�2s��̕i��+}�����A��E$=�P����������M)�Γ���xu�y�D�N�#8��͹�0�@�O;�ߣ_��V���$�A��+����*3혧�쵦�}8�'�W���_��9l���U]N����a�)*(�`����@+�����׍�} �@��M}�ͱ%
��S�����W��.N��4�1YB/��vP�N��[������ޠ+TqG��
f���谰fP�ll�n=^���4n�,/��	X`V
�e�{du�+��NsZ#F�>"gr0 %�&T��T`Ӥ5�|� �/���ϡ��/Q�r��Ή ��7=�Z)�}��.�C$�	��z ����-A����\mz|/z��{�9SZh*����Lڞ�q�iA��S���YH�H�b�!�a�IH#������Tp�09=�	�h@r0�=L]%nNbZL�#w���l�)�S����H޿ؒ��d���m@r�"hw�i�)�̋�2Yo��jk@�{`�������1<�L��l��$H�nT�vM\���y�My�Ie�@H0��Vҭ\�k'H�yOTF�#A�W22�խO���w�e��(9�Rn�@ꌧi���!=$��f"�7�@�!�5�4�8\��ԭ�a��f�f��ee1W�߭��>�܄Fo�q����|�TY�+�*"}d>��Fms��f�Oa��B�����%M�t~�ޭ���8Hkl:EM+
�+JÝq_M���d�-0"�M/�ؔj�[���VCb�h꥿�z)���l.�}��<�G�H޲}?�f;}�+�⥥s�W�y�h--�����ZF�(�~���?�n������Џ,"o?�Jk��,UZ�x��v��茍�U�N�k����s� -�Wօ��.;��Ӓ�J(TO�����n׈j7+Ò��o�;�`��h�5ګ|F��@ui�f"��lي��*����]��>��-��y�Wfq�㛆/�#*E���xN$f��d�����ׅ��
Jj���_gV�5ԕ���
��֕�땪�x��������b��i�)dyG����u���v>�Z��<!�)��_���Kߴ�����^��n;$%*^c�2B/���,=�����8Xq:][1����/��H=���:�|_M�����	r�b�4��"�����	(T�&N8p6&&�gE)\>��6���L�D����]���blC�y����g�A5�4�d���%0�2Z�Ӿ�ʪ(ڀ܁Iե���=�A$�u�5��	�M�}Q�d����NY������B�-���׻����X�j��a���)P��뿇�&)Eˑ�i��an���+�Mx9��tN�M�H'�0���WJ�9���vBt��!����u���6#,��G
�j�\�vm��@LU����r�sq��ߵ�;*�cb~K2�������9mgg7�������ű«�yLxKFW���ƞ�K~G\�dl�g���]\Ssa�3ɿ�ߨ��+p�LX��|�~���(���j�k��-�Y:i/Nz\O2��Х��}�7��V�.�����zX�3�LF-�^9�ir_������2�4�,�f�U�4�ǩ����ScI�i��y@����Q��NHvNN$�Ʀ�Q;��F
��6�b2/�,]}��O)|6�C��>���$"o;[.*�I���Q��4�t�b�q:d�&�PE
�Ν��(�<���2�nrfܾzu_�������	�J&�+G(7B���I l^>�{xG�r���"v�]��&?���v��U��S�J�+�X�^��d�Y��X���ȌQ��7�������[��Yvw�`}}:��,�v|�8R��ق�%[�h��:ٝF�_]�~6;y�١l���i{�N���A��޽
-َQ1�%7�8V80`r�R �nC�ve)_\��K>>��F�:��S�M��
y2���koW}J7$�<m����A^�ʥ��.����=�w��.+�bUC��}�I��f��� �`�8X,��hF&��h�#�������2U9G��YlK)���^�#RR��K�E���	/������1��/����r�7�>�EP��&�R7x@�p���ano/�s�xj�#CYF�t�f�zc�жc�*"�[�B�x	��1E�¶dIH2��Jn;_1]O�<�5W�C�=��G_�
d,{���Sڬ���-��mX�K޴iSI��0�n��{����
�TE�b|���"?��0�����|�	w�g�.�F#V��&�>��l'{�7[�]9m�Y ��%����[�6��Qr����,��2�DZ���\�����_<F=����y��۴�=(b��Vbx�F��[u�����H��\�c�=1�@{>�@_��aJ�'��!U��q8�al�ȑqz��W
s�v) J��9�=��~@Ѩ�~��N�p�v�)6�}T��f|'����`�*:��R25c��>2�&C��*za�`'$�̟�v�Ŭ�����A���.��,,�䣞�3�M|ؠ����	w[�W�}����
�B���a�"���`#�S��Ĭ�ج�;��£���0X�^�HiYq�ۄ�g�e�c�TI��
�4�M�+s�M���8IZϨ�PDr��ў�����K�w��d���Ҽ P�)%�\)���!��/**�^��}$�>/���G��;�l�v�˶SW�6�������D�w?�Ea�r"��u�K���v,e�HD�:E�tݤ���]Y�M��.�R�,�t��'�����n�|����^$e)N�E,�{��8���-_����;?-�4��߮�q�f��%��ڳa�%$Z�Flww���5H.1m��{�r��I�!l��;w���7�;���0L���O��k����9Ӟ��053#���<�)xLBb����:�) �)^��7���{��г���Ff��8&d�%�3݋Ǹ�n���$��I,���k�a�E��(��-X0��=�g�s@��8u.�����n-����z�Ny����� ��޹��G�AR�)e���r`�ᙃ��r�>J$������CO��B���~��Y�|3B�7'��t��1U�����54�pqq��� ���OOPaxA�t�ڳd^ }}�x�6�5�L��� �'&n�F�hfE
�� ����<��H���>5>&��hE���4���Uss����j�'�c̋�.0�ќ����L��B��;��<q�̈́q�d}0&B)��<h�ƍ���@�Ѫ���e��6�! #�w+&|�1J�9ި��/���Y!xF�X&(qp+P�,l������"bV�
I|h�)��ՍQ&A�e�V5�T�X�c-��f�g.�O�����F|�!!��@�xf��4�����Q��7�2��s,{��f�>�pbeeg�:������a������
��NzT���Z���x���@���-��2��}^���]�h󪲅��\�֡�1o�V@�7qq���uј$B1���d~��
~�F��y��#;[��x_|��j�hw��v�+Gl�Ϟ��k'@�� L_�a���.�I��)�l�w#Âa�c�O���8��-7X-�g.�BCp���nX8#{�9� ���HE�ջ�28!zޖF�{::\��+c�������h��ڪgnn�]E=ѹ<��S{�S!~�VLW�7��$�,��s�wtt�����\�c��{h4MVz�\�=s����6p�݇��===_à�����Փ��)���M4'��i%d�t�D�tyQ��d ���Ъ�<7�!�H��*�1D�6!M�d�ک����=@Y�e"|�#{����۱?�5��-���T�R���|��cf~aA�g�祀��y�> K�I��¾>&���#���jl�UE�h17O���vWtt�	3y���C����;x� V�H�G�Gr�����[G��J�op�m;�a�g��ҬR��=;����8��B#�@�c��1�o�n+�+҈u��7�b��8�SH�*k�WN�G�����d�q�����14Wֱ��lM�Vɢ��˄�S�a?�]����>�촶�����*)I�F�6��fؼ�4�hn��N���}�\+QT5��?�:�6��t�Tm�D�F>�v�3$d�m�V�fb��<1-M�gv����]��������JryW�:hh��x�UtG�?A�"���3����p�6��\h >ؒ��y7�j� %�)ioz���6�i��K���+�c��Qe|B!�bء����*����Փ��B�Wh�N����K�������'0ݍ�6��L��?N7m$P@�1&��%�'�FT�(��	:M�?��2���U���}�����k��� ?%����U�ꂉ�����������*TcҰ�R�/J�\��#pB�1U"*v'��T��H;~������-����0����=@}	��
ВA���>����=�F`rF���1�E�|(�SE��m�@����6�C�rtrR3vV
��|��sW�;lX�|�	_Aֈ]�3��i��?b���q!t/��[�����m�xs<�B@o������zu剷�� ��u?�Z�L��[����?E�����"f9f	�����A�8W5���>�jH�޼���y��h��OW����P{^��$�"�:����X�p�`Oqo\����`dQ�Ճ����C��6I-'�bd�-?T�e$���##����Kg�b�iy��چ���|.�!�m �ސ�wF���{DpP��q�%)��V^�́ժo��XҚ���:��.���w,�#A�<� ��9 G҈U
�G���8�0F�{d�i�6��J�0@^<�>�O�LA�# 6�����=�U��r�?��Z�?�`c*\�fFR��v�A%����� ���zК�;6��?.���ۢMS�(3c��%� �*��-F[�)���g�hy�f3��Խ�6}`x��/��:lO����Q/���n�w��bn2|��2�W�1��*�V&�Tَ4�Z&�SB�!x�{��E���b.\�t��r�;�%�N���m�����A�'T,��$hhG�=�y�hܔ�]��������rG�ٌh�_J���^����.���ܙ3�Z|�Fb՟ _>-`<�٘YY+:y�鍓�'_^0�j<h�H�[0{���~?m��7�g��I,ި���������I���n<5��1�����2�.ށ]��_�����
b�,^D�>tE��X�,�8����3�����Zئ�_jeq��4]ᤠ/��C0����2釉�;���V҆�R)�]� ���0)�d`�i?dsO2_������)E)�NI0w�%Q#]'�|�`�	��Yc�j���eה;�3I#���e$��r<���x�&KW)��Y�Wa�+��B	�;<+vF&B9�n��'ɽ���&���{ϕD/�����L()�hG�3;SE�RXx�WY�P��k�g �M���\(/	N�W@�`k�2xz�{�&���=	z{>{�Ī���x3]�DnS�5��4�VQ��R�m@ං،T�����4�`L�&���{���i{��S_��a�W/1�O�]�`o�w��Gц�ڒnj�+�D8HX��'f|�v�'jj��>p�5X�M��� ��|U]�B��K�6rG��b���F�0�#""\Y@�HU�����9�W2�\[��)���1�W�����梩f�ٙ��D��¨����m�)�����
�Qs��+n�זC2���������.?�aw�B�:����L��6,��w������x�VS�O�C���YԺ�=f���[00(�~Orr�2K����L��X��{�K�
���cOR�-����� * �֭�4�t\&�]�� ⛅O�
�ذx�4��f�(�߹uk-D��)���� 8x���͛K�*C$]�ª�u��}qNN�L*ku�\6�fJ�#��=(5����Z~���WBq�����/_qv���d�y4i�RD�Wp�c^�R[�T��U�q���ۏ�F��	Fb��ѣ�\gÊ ~������7.'�~~��3�1Ug� BQ�n�/�i�_`�9�O�I�[q�yR�~���H2tv��/��	�e(.��E�6�!���Pr�L���,���v��s�;]�b��z��0[�G՚��U��z�?=d��-#����\�2)2?�N���ÍIxM��s��son�[��a`�c�ð֧�2/�L�����7zA�Z?l�+H[�vv1U��۳m��W`�'o9v�ϝi1%0�k��F�b��zϟd�qzg�N҅�{aU���LR�`�`���7@��T���M����.��'D<yUR��o>�=�Em��?rL(�L4x~bo���(w�����6r�N���I�NEr�B��8m���<%��[��'��p�Iw�/Y'7P�%�������x�e����f��Sw�и������;��Mu����X����Ζ^�l���t�ȕ�����3ݎ����,��R��^GȪ��n݊�/`104�_��k2�Kx���8�n$%)|�Þ*���m-�"�zX�R����.�	�Ô�2��u]����v=!�`0������ß�c�l��,K��i����"�+��vc�I��\�4P�:3SϨ�ÞH�L,������"r:J�8_�Wd"tfEF>�L����� ����p�����$Yq����$V
�C���2 XՄ�)�t?)1���B�B�b��l?qq�7��V�>w1���n3O7�W��@x� 嶤-Ex�*��\������[&��7� xE�8D��G,�h~ZNP��M�SB����Y������� jO�QbN�e-���H������ `%��`��8��d�3$!����}*A��;@�G�l%\�.؄k�􉲜�<^?W(~�
�m.��<[�	��i|a�.S6nKӤ^�T!KכvڢQ��YM��a�y��/���$���������6r�b6�7f�Bv�'��í|����v��A�h�e��š��4֍nÌQ���K��G��,�Pc� ���ާ�Aߪ�����`>��q��"�Y�� $�ԩSy��||"�rHp��vb�@`�1-�����|����ĭݟ �xR;��c����^����;X]�����%��D��
�MF$mdl��~B�L>��&����&��0H�a�)<
���O�W��׫�5��*t�=? @��yk�E_���욨�+�q�uu~i/!��&�}K�`��m��ok���iʴ0*�΅����{�f��07��J��w7[�t�C?����,lYdAp�s��I�ֹM�F	�
,|����=������6���.�2���5y]�֮X��Tj&�d���*��:,�ȏ�9<����%u�.j�]�v�e����a�g��5m�N������jٖb��_�� ���:�2�=��@\"���g���KՔ��%��|}�fh�?FÂH��'\#'P��4IF��?Q��ٵK���<��)t��SXTTt��<��6[������2��a������ק�] SB����a��A.)z�9�p���Czk��X5���R�:����Ae�]���7p���
g��a^���C�����7�?�J���_��K]�W��G$��t�6ƪ��C���槭xpU�4�ʻ_g��ϱ./u�Hs�w�{M�����ux Q+��Ex
�2)�u	H8� S�
�t�/�7(_�����SkQ&8�Ç�Y�\+K�Sj��d9~u��\�q��VG�8ѕ��sr��ج����֔��\kJ B��
%�ӌħ��u��[�-MF>%v�y��^�ڗ�<?�4Bb�c�����aEz�Ios�t<:4-7�_lҮ����!��Mf�?��_;<Jp��R����x�w5��/��{� h0 �AJܙ�C�H�%����"�y��$� "�òt��FO�q����� �:��(�����<����]�W��>��.�LSK�,�|�o�����9�M� ��<��*g�N6Z��.���	����ծ�|�f�/�{�t�X��?��6»���Z�.�w���tϮ�.��Uu�����66�%� �Dn5�3��tU{�g�T�{2�D�E�2y��؅m��MN?u�����Q�U��<���c1{-�]]�!��t�zuz�U�<�5V�������R3NLL$M�"i˙!�ś��2K�� 9 v̆�u�r/�zI=H��u1��͕�0�т,���i�������b,�$*W��=�@� �O ���q�ͷ_�
�I�8o�z�VK�!�/М�S33���0�od&ӜMZ�AfھZ�G�lW�5��ķɥ;��V_"�v�͆��z�~ٹf�,�}#����ov�WZ�nd����a�������Ӊ/����������arP���,Tc l�tf����`�r�4ʋ��QO�ż��b���>H�6>->���C@j���,��e�}))�������o�myt��~�$dvq��^KP�L�'�ج�m�W��b�p�O���Y6��NҪ�-5���G��NM'����j�J��J{z���%6��r|�r[����f�����Aڡ�,���f�C|�y�w���/o����޼sl+�L�� *^�n���2��%K��)R#�4���2X6��֏�}9ߤ����+x�2.�abZ�,`@��4T/V���%]c(a��7<a�f�邚ȶ�S�XRK�QG��a(�3�MX�)S�č�:qi�
�����R�v�ik��rt5�*��'��v��aǘ�.�]�/ΑNL�C���:����[ Ɂ�sa������>а�5��0׈�/�*֫��M^|(\?QH�P�`����Ç���R&OA�cͰe�5G܁}�eD�C)�#6�o��`T����l�����y����@�!����x�ei�5��v�lW.����
���	WApG!�i֦v��������L�"���6��Q��ӳ?�-�Gn,22RE P͸�PӲ�eݲdH�K*"���c�����C�E�v ݸ; ��]�[��?�~�R���nA��OҴ� �q?"�thy�s�dn���E	iF�hrrz�2KM0:�@KeW�3���3LȚƋ����?.V�Bp�x�315WE���3r�\��c�/z�~>`F��ggٽ0��[��N`���S��P��ʂh��>��?ءw�(Z��h0���)Y�399�{^hrE�������%��"�������ץ����٬gGy����j���]Җ%&�	K��MCq�ef?F�c��_�빟<�4�����o�0!k��վ�2�7��2�s��`��?^�J5Vx��J�c��Y��lI ����	=�@��e��!���o>*C�<r��?�h�-Ja>r7ֱr��������S��vE�m�h��9w�)�{��]��_ʿ��߶la.׬��#�UbXG<_���d7�h[��y��7����$�rcQ�3���J�q�d��:8k��n�Fe�� o>Q1�HTR����z��ʪTzeeէ�Ƙ�߀_����b3H"�yg<	�N�%i�Ƶ����A
��lŚ�z�"ۑn��{����~��Ƃ�*1L�򆽎�h��YDx`��Y�^ܴy��#X����w�B����ğ��mt�R~�r�����+��y\����j-�#��oE�q�yze<�q�&��DJu�Ԙ��� &y�R�,f1x�4"��s���29vb-2u�ϗ�kע�'9�v�vt�]���G#v����4����	�;+�Ԟ"�_x��={��H�c�^��Xﾚ�D�ۀsC����>BySS�=5|7��Q7�R�����i@�'+ӳ.�g�-�BWE�ZѲ~�,�9�ng���=:\�2�;!3$k'ç��ꂠ9�Ֆ�硝�툛~~H��kݧr3f�u�8���^���jO�{-��o��v���@V���C�&d7���m�]����ɑ��Wó/����qi����W��d�nza>B+�e9��lm�bz@�;��o/*\����RO{� �*���"�y;�HY��t�I�mq��T"�K��t�,�:Zl�dd\�ZZ�@�:���콵��$t$X�_Cҫv[�$͝��@@��"���U��`������odM^(n�V|hx�j3�@E
���Z�IiF��U?l�{m�j<����+�~0s>&���q�R�yk����P'D����Wc��7~��⪅`I��ɧ�6��'NDG`��>���%NNe�8$`�x�$˗��� �Ng�ö���px�4GG�վh󪘪{�a�xyy9:���t�����^��O��_B] ��7��#|��B��˿�W���2-�����i�31�0s����T��(��u/p�`	3�G�[�Ҙ]����`/��o	:���	��Ǉ����rz=�N��N`n�P����j��x��\��ҵ{u�W\��މ/����v��� ITh���C��� �1[Y��)|xϞ����p?�J��d�G�n��&��mYV���7�8�B��l��4���T;0�����~�ؚ�Tx3lV(u�?4!����f����V����
?�=@���;u��e��ؑR���yٌ�kƶʍ9m8_a1�A�ѳ����s�� �Y���9ݤ��6�f�T�d������a1����Ax_�����^�i/ͻ��s��3���@`
f]�Y^���q3������s�~f�����8���ǹ^:��_k֮7is��sj�)�|�mq���Mw������ռ�}Z�@<1.��fz����i���^D�����R���rN�Ä<�[�M8��f@��_���d�� ��t��ޮ(�����_���_#R�O[?mgcS200�_p4�ʺ���m-)`���D����0̰3���i�F$�uUXn4pk�$3'}�	w�}���bڬ��rcmO�'{ܖ\��Fg� 5�X�P��?�l9�FUj�Ȟ1;=M*�Q��$:j�QUA����x,�mH�~�+ى���сr{'@%	*���	�zp X-@�8����C�nq���#Z�����C�R~�L:
��:W�ֱ5�����c�3�?��^A�1�v�x:��x�E�r���	F5��X�.�����8��'ؓ#F�qc+�'�" *� ��T��~�V�<f-'�:�7(]Y6qsv�Gs�N.ߠFq�`ǆ�y�6_	��c��9]�D�ښ��{�Z4��Ar\1����M��ã�6~��l]���uia��l4т����9�]v��=�ѕ�7�k�A��JQtJ���|ie�����l��ů�ܾP���D=^�D���,]o�dQ����)+��řV�?��[p�hZ���o���Kc�Q�@�}��Y��P�����FU
��h�2���xg.ʄ�p�R�� ���gNoA���+�����g[J��4rB?���X�Nf����Q��7vyɱ���,-����-�q���e��:������xX%q�;:XCfaayT��+x[zYĲ_��J���,c�t���1��]�(W��} ꖜ�Y60`�V�ø�:"�T��Q_H�o�N@�����iǡP�hX���X�Uk�AG�<���V\iC��+�kp���)+�z@ب���e�X�^yNN�!����[�WZ� �)s�ssW�e<W��&���,l �ucc�t��-ȭt�����U �.�g]w��e�Z%�G�l�IN"W{w���jQ�xL6*���P�|w��y,�~�L��Az���zÇ�lj'\��;v��m0&�%&&1
.�t0v�ZRE�]�䴶��6Ņ]llؒ��׀W��p�[a�=�l�y�Ȯ��X�|8}��@^�*�z��ږ��
sW�9a��̉I�����1!��%i���� �ϰ��1�4ܯ�V�h�����8��ݕ��Z�\$i�����a���缼pزߠ�<p�N��g��<pK��{��s���x����E[g3o�Azz�pS�
ox��\��[��Z���}5�w)�&���=���9������ޫ	x_�^�>Ӹ\��$��߻A؝�j�����k�I�Z�mڷp������]㛛{�������ݗ����;�R��~^���/����&�e��z��Go����(�Cڕ���4�d���+�m"�����B�Q��c^|���J��׻���BB�`�����ɰ񁮢�\��A�/�;v�<�å�������sp'{��%i�����tZt4������?8�Pe���>lQ��l�樯�M����&�?��'L�g��Nxz$��fUد��z�Å�A�q��ә]
 _i;��ׂb��r�&/O����g���K����9U[�j,8���Y?6�ћ���H�E�]s��=x��eJ�ȧjr�-AF��i��˯�s3Z��߹�ٿU��9��)w	a�-Z��ˉS֔�i��y��x���V�wG��G���b&=n���j*o�tPTT�Z���J�w<G�w�aL��s=�A����}�Z�2d����ǞkE�d�W}���_�ҡX�	E����t~�K����#���*akN^ay ��i��O՟����q���w�|�n�ڷ�3&?�p��3L�M?O_pD��ʥ�nJ&H�b�9J�ܥ;��'$�Zw<�}������c�~��s����Lѝ~o�����=���c;85X��Ln��d�o�a5�G̛�q`��`\�������ԥ84sڿ]>���汗Ns�]ͻL�U�/)Ӑ��1&_Y���}�(���#nǦ�=;�+�X�_�pџ�?��K����O��8���w�w>xI�v����I 5Xܟ�.N덜�b:{U/�o��9ⰵ?���>�{�A���9N=���B
L)�Ռ^3���wa��gnf�5(N��v���-O�s�x�=hI7�rf纏����W?j�0>������/e��-za:�b����{�k��������5ΘG��5ȍ��l�vy�V�7��1&�_���j\'P�����
;S?�m�k�gbb��4pu�{�����8u�FF\#bMk�Ӵ����7H�H���J��@���٤������`���|Ϟr?��̣�����-u���g8�K�D�]A��#v��_Ue���+��y8y�,�k��f��l������o9[2��%EWռ�7d�j���d�CSk��w�9̤�OoR�]���\dpD�C�tD�p	����_�s��I��kM�7lؐ�8�6��z��܇I)�G�v[F�O�2;�����*a����g��fh�!����p�'�r�˧W}�UH��>�rwE��cU���6?����0��qk݃+�Zo5�ut6HV��L�n�������Mo9�x���1��^��?dF��ҽ$ey�I�i~������G�!p����zS��)KO?��*��/c6��� {�y2F)LU$�Ar<7���� ������٤;����8��<=�����w��eFe���[�Ԩ���M߶�%K��(o����7}�?Wi����Y�����3�b��W�W�d��9mC_�UT+1�}*9�奤l���'1���Й���aw��g��x�x+h�5��uKD�nc��$��W+�z���K;N����r��
�g��A���D��-��k�v&q�m�-Uˈ-=�Ƨ泵�,cy����>x�-���~:���yzp:%{����gk	韖N�j+
��=��b#O��*��𒳡N\��w�4j+9"vҸ�=����uG��;"��/�V[['���	�&I����s��ǫ��6���`lM���zIQY�g�3�iv(�?��u��˻�i��.�R@���oUcM\\��9�������C�*:�����a�+��z�Z��G]���(�LO�tsVAd�id��L������)σΪ>���O�ˣ/��>����
�L�����=��e����ۼ�,3;�j� �?{Eo3S�p�F����7v����o�Iφ�-=����/������4ڜj��0�.�6�����R���p��}	z�jit��_��$ ����!Y�������`~P�m<�2c���8�$�k����x�n	Q��޼3YKA�Z� �����\�յ�~����t���<mӮ�<�9���7�x�ݹ�7^j�F����|Pz�9��{�ii�+��T���:��>���r����t�qю��M���A��בg|�s/p��!I�Y�G=~>>��'���&��g���Zh#��\�`LؽyE�VU	��SJ/�r�@k۬7���v���&''S�L�cZ¢������;�ͫ<�*˃�lb/�b"�1
�4�����=�I��= 䊨����,��ߨn�D_������p,����T�$IFG�
��le�gvvFh����l/�+�!!��MIVFF����}_�����s=׹N�����s>�w<F8DM�b���~<s�%��������Č쨳�S_S����"֓ٓD/����<7	��<����Q
m����hC�=�K�~\K� Q��7=e��{:����*-#�iA~���}F���hD~6Z����>��IG�:�������/�����b�2�ѽmQPD$�������@g�@�ӹI� [+Oi��L�� <��L�zg��S)ޫ�G��=��o�����ks��T����Mon�0{s���-���Or��h�X����:������r��N�_�
F�sTA�9^%���f�	�슌���zeBu����������{�K���oԉ�B��=��H�.O1F��`��Vj��~G��T_OQ����/�[(�NVp�b���+�MO�w�/<�Yj��C��Z�����b��ϓ��n�.r�"��"�_�$�IJb[����߅�����Ӑ(\��9�vs��P=����oԅ��F�B�kK�n��L�P]Q����>�}��R7�
JK �x��?=%/��V9p�'�q7z�ɉ D��Wo�{���B�}�6!1�B����)��|���)������mm7��4�Oy���5�T7��`?��8z�<T.^�(�}`>�m�sm�.^�"���_�!��gzĚo`b��־_��Z�������c����Vy�-)kG0�x��,��fa�#��	�iߕwB5~���^�Q��-�8����s��P���S�"��c���5���Nc˗��6���q�}�����pl����9�i�����n�����h�b�2~��'u�Lt���@�h��q��06��Y�H��R�zg&�*����)��1��)���	��o�OIVqfLN�%���v͛�{�g�����i>~���"�{��彩A�נB3��5���k?��sO����f �L�����I�����kP��U���������U� �Ag F��C�k�]���M��������s?�kfr@�:3_L��W�'�q�B���`T�@gg�6ɕ�J���G�D��3I�-^I}}�?�����
��jL�Ŀ|��#ÒjR�i��؜a����z����/7�gU�6��s�,�s*Y��Y�<��:E��W��P���{�����賓�����߬�!p�C$Q�nN�W�j��Y����aGʫ�ˣw����{��FMvq����Xx�E;!G�^A9�p�<�_�mp0�������''�B��|��!R�eN���}u��_	2�Z�p7Qx:1^t������f�&A���,q�ש4ҹta�%����p:����߮��<�
qz����bu퍊�D������Qξ���݇�޼��*��K����#��:$�O~{�ܽ�@��!�ԏ8hC�������{F��L���Ui��k6�rZ�7BЉOc˶|=e]��Cc�6/�D�H��{��s��S�vΏ��~*ė�*�����.����aA ��C|\��Q1|��9K�e
ܙ[�2<-[O������=�BK�����^*,g�;��;�`�����T��cK�<�Q���D1��t'vxH�߯��j6Zhw�`�6�-��P(���K��\?�.�����{�K��4<�Ć�,36�}6�����2'���y����������|q�}�&�ϼ�ӦW��Ry��lB���)�	��p�4I��/�c��g�M.���&k�(�?(N����isy���Ə"Zn!��{���:��Ӹ�����yj�P]`]r��O����$^B��+�A�C�,�iѨ�o�y9�$5L��#�	���zc���_��`�����_�ec��W/��1�`�>����$�`������:�
O^�SG���������f��L_�����f�4��H%v����/����D�|�F��k�89S��N�1��]5��:m��!w~6�_ ���q���2�MW]M9LxAQK���l�0G�J7Y�I�~]=��CJ���p�������Rm�D'YG��q�YT������6'7�!��f�Kh_T��]M��|{�o8����EMI
=�����_����_�4~?�@y�%lowp�c޸��S�F;���=�g���z����m�����w_k�jre �rӆ�̷KX�.�Mod�s�r'�� %ѻNb^���0\Z�.p������en�=AnR�lC<	߶���x��LJKο*!� 1#�U��M�cHW�9q~��qΔ����Զ͡��L�󝕄7U�'2N������Iݺ�"B��(�Hcؐ�cI�}�R\�C���f�{��t���
\�?��ü��;��P_��QL��X�{�ɵ��j�i D��,�[�/d��hO��9(���؟}(Â�?���uʸh����N�r��a�����'�����sE�ox�:�[��5��Kr���i;��;��;�)��w��G��	�~U{��9?�Sx��v-Ƿ*�p�+ �0!�1��묐?������]��ݿ�xl���G�|��bhl���Im��� :,�q���$���_�o�
��4ϝ;�,�9�O�0�JjN</|�^ۄ�\.��:�ȥY�B��h�L{�����1xE\.ؠ��k,c^�������V�7�^o�/���$�{��}�sR?�h��*�����Y�<��\��d�5֗����7S�>�ct������m#��W'P�p�����z���TI�"~$�C��~�3>|t"�6Y=U�nʈ�c�`�h����@j_��,���`\���X� ����c��qζ���'Z���6�A����d�6�o�=˶����&Pz�,Y�⟠�����P���Sh%*ɥ�Kr��[�xب,�J*̚�����������9h������v#�<�%B@�{��鹶	%�?yT4!%E���T�h�V� M�J8�>һs;3��I	י��鱵�t�]���ӿ�%��cup}}��Νݩ��_|�!w�����"sߌ�{����'t�8=�;�a����h@�)bzi��u5���J/yT��C��A��8�!G�Z&�*��<���7�Hdй���i������O�l�����'�ۯ���}�;y�Vi�M�b��fT@Eo�Mz�+�d]�v��d'��<��|�&�����W�v��W�Q�TU�{=W��<��ɦ͚9A"�X >����neg}_�{Z�]�'��e�0�#�^�r�#:>TS�co<(Uy�QP5�c;eX��,�B����=Ē��0	��P���9��Sd��_Zڨ(\�W~HR������K=�CRW'9g�(;ز�5���^*�[X�*h��Ə���lm$܍��ƅ����w��8��q*?I�bf#��
R6����ŕVT�XW>Oq5^I~=FA�v���CGnj�,��[���-���8
W�a^�F}/��z�MT�d��㕸�Z����OD�3����K�LF,N�9�
(t�o�'���Maˇ��-n�D�	�k�.�G�Ug_m`/>��v�)I:�$E�Qfއ;͆3�10ɝv���NZ&ݬb�QQ�i��i�d�S�{�	��&
'���ړX���@�J��U6��u:!�VYy1�����
���֥�q��|���o7�.�R���㶍�����p�T�St��Cn.����ȇ6���Ʉ����\��WJ� ��^�*)��e�����jGЕ�@��G�3N��{"��ݸ��ݟko>��|%�jw\��a26���l�7�s�J�6�]U(6Yi�:zݐ��/[ƺ�V��m��$�_P�NR�+���1$����~��8K}@��(���L�=�:Ÿ�FE��o��:��u��WD�B\�I�/1p�P��ipSnu��u#����Z�d�Fvj���ŵY�:�N�y�uG��|�j��=B>����$�mk��D��V�� ��[���4�;��'�h����#�� x����.̼��K�]U@#����vR*��.""R�RT�H]69%�5���$y`ʯ�����G%���^�/�7��rȰ��q҇�;99�:�^�e
�<{�ӱ5=��|T�%�p�`F*�ϩ��5�_�ܴu���!K�x��N�����L�Az�f	�n������_��o<d�&��[�y-�455˥qцN��>=��J&?�=���*>���+/+����-�3c��&�֪����s��E�v��l?3�k�PH׸o������(��c������z�C�$1ϩ�|�����2һ׼��{�4X�cu�A�ʜ�[v�:黎�mVn(��u40������H�uu�)㹄�� ��}.s�j�L���J-v{���ч����:y��os��-R��>ny�v͟>�*�U�ua�6G'7lYg���N��hP�]H�uU�v3�_	?���~L�k-zeU�A��ӽD�;3��"���	�*�	P\���x�pQ��f=��I=�mY����$qo��Ռ�̀��Y�n<���z�sdt"��dUԦbo��N�v�	^���&^o*6�ލ1�^�-����m_�����q�%-vzj?���j��ێ��IM13�_�u���s�-|uyhS������������F{8���Ƥ<�������=�?cވ>��yû�;m`m�u�qi�/���#Aq��kV����j��g\��7�ϱ��'2,GQ[gm����u�֓��2��x3�x2�ʆ���-�7n��AJ�%n�Qr&�ۑ������}/��Ctr<���K���/=E�V���?o�<�u���V���O�I����w�����E��ͼ���̕��=�� rvlل���蜦{6
�*_���]��ݳ�ؠ����I̸�����m$\8�~���&��e�Q�r�N�DҞp�-.u(�M�n��I�	��ڢ��`�ݜ�y�l$m��-�3�!�7ؿM�B�|vݎ��faeL����w/6���pr2.e7�۵������h쉼&sV5YH�b���X���K��#A������+b���;�(��!����n��Ι��:�7��&(�վ����%��îD����t��b�0)�t!�&mllB�k�g-����	�h;ym"=Τc}���{���bC��کjj�F:Ž�A�/��]b��Z�_պ족��D!'�s�U�L6�D��Pu���C��T
��d�K�/���:��������DH� ���5i't�f�4�
j�_�8_�L�9��Dr����L�b�~�'�z�)
���X�ʪ|���^�K����ָ52*��)	���0RڄN�ٻ
b�϶-��y����:���+N09m׌29�Pc����D���H�Wzhg�Wz�_�3�d%w���Ҫ!5��W���o����T�.�g�jRn[�PE�.t����iY���K^j�Ƅ7����s��� |岃��MTM��N�r\RU,�Bq
��IZ\����1ڪZ9.7J�R�J=�O>����這�C�4 �1���	�	�������:�Ie� �#�%�s�b�??�D(��h݌u�5(p��}���OYaQ��)
\5�'�0=�kd�1a:ame%.7��1�V(��Ԅ��P��j/���0eL��s$�Q�'x�@�|&-N������E�?ST� K�BKo��_��Q��ڐ����P����٭&A����{|(����5�m|�j6�'`X#�����>%V�CR��'�;��fAg@�p��t��ri�
�ͮ�^~���������IҒ���ȕzK�L@g�u��&;}���).|�ϑ�	%eeΨ�O��:;n���?%�2���,��&�m�)�7��R���D��"�}�4�QH/�"�p��+�x��6���}.��
&ٳ�������7L��Պq��i���˜@��$�g_�����L�M[GOq�	m�{����,4s���*Kb�o��/�(%�/-o����C/6�����ͪl��*�@7��dt���(���V��S�a�G^�Hlm.�Snm_������O 8f���[�����:ۿ��S��|��궷�b?D5��:�[�+�(���-��P�C���U��i��恱��E�~���Kl�)h���Ռ	��q��s�%?��R�2F�("�X�$����+�m�	 �+���L<:��uks}�xK���8�3���e/��ۅ|@WkS�i��Xp2$5[O+�����g�U{e�2��?���&3��)�I�h�du��]E^��'yau#��ln��he\S�#��<Ċf���7����'gʇuꆩ�;�57X�c��zM�,����:���V�S/ֆ��u�+Æ:���`�s̑=w�f¹�b 
���{�k�AH���	�4Y	
	�f_����<�vUa��'�����`
ϟ�O"�����Q0�v�6�� �8 �����u��*�!��ԝGQ�D�������.��Vsf���x�+,c����L�m�`��]Xm�]~���<��ْlP�S���T����EM(�j%r��9]Brr����/�#~9�{D8��U��0�*��l ���������I�JA�A.�YNql-�ې�������??\��i%pRr�W����"��PS�10�,9U�2�3�Z8���F���#,\�||ƼǾD.��N�ۃ��
>�ɹJ�J�pZ<\���(:�x�ȍ4�6�W���u4#^N�+2��.0�����\�-��+�l<E���$���c�ȇO|M��;�[RTD��\�ͽ��)�$
���t���O�K�c�Vs(���!���7π��7x���{��onڔ��46<��T]w¹��eEd�x���9Ӆ ��� ��yⓟ�����X����K^�ڼ�_���`q~x�r H���0�[���2�n*�|Մ�e�8c� Gm�Q��|ǃ&��Vd��w싱r��3>Q���}����͉<��9J��d?J�̛�A�,�ϔ/�����1�Ӛ.$#3s�'Y!�)�ZFb��2g���u�pa��ӛ������EW9��.�����.��v�e��K`�y2��}}}5�����T��7�W�HQ��j��@�3‧����i��� ����
~�����:��8���x�����9.VS<�~&|j����f��.�ȭ�L#޳�����$�ʮ�K�H� R��p ��we����Z����Rkgj6��O��~;��s$��,J�h����8J&���5滨��Y�§����]��Y�1�1�3����p鯿�Zq���KIu��^q��S��&�%�nLHH��>�?�ArQ�!R57�Q2���M��Pu��w='��x겇 ��a�������`��6� ��7d�ڄ���!��aZ�)u��jA�=��$$�'&�����@�&2mK��h�0��P��Hm��[�H9쵃��N�;e�ϡ����7k��`��!�r�w�D`�S�S��Ԟ�������a�d]����eLXYp��D��P����4L_�
 <÷:MJ��\v�nqE��1�Ǎ�ޒ�hfWb�	K䧝���t9�ʏnen�)��L�R' ��;����;�]Cè9���H��SKk9B�k��ݺ��|c쉰O�b,�ߝ��8�z�2����+�I�U{��M��\���)/S�ou6mU��:���¼�a��n-pR?�Sy�
GJ�Ebd��ZA��&R,�������Q��ĵ�/�
R�s����+ks)��/���:�?�Ҭ:^x3�S�<o�A�C��2��������{V�{�M-��4[����u_L9�qq7Ƒ3|�'m�`�2�}]賓%~�Xru	��>�9%�y* )A���������ǐ�1���]#)tk���>CU}���~�Q�x����b�5����2����3��o��5���J���g���ůt1Rt�,�l�1gᙳp��:u��?�)�[w e7�W����hjjB:(/�Q\���� 57�KjP�?�yb$��ai\q�r���̝(�<���� ������#Z�e���Mf�Oc�@���<��� ��ϕف�ԏ�l�R�(;?��k�۶�Q��!�b,'N��^�|m�?��S6���T�������b���0U'#�� �#�no����_�G��iUM�Zm��ˋ�9���VC��4u���i����lQב�����L^�Sg�k�V����լ,��m����E<p�E��e_ӺT:?=P��~m_B�L��W9�<is�+U�Z�<v�L��dʰӞ�q�c"���Zw��5P�w=�z����:�����w7	hF���~<D`�dChh�yc�S�4�N�(�u����,&��{�v��Ё��'�n�esi�8���� ��Q�|ß3q��$���a��B4�	 HG��O���ku��:^j��K�,��i���m�����AZ�����W�1�4�/e���6��S�|��}A*�6��ތMq�B�K�ē����z:>�l�d�"�zV幚T
�e1R��������l��S.���\ް(Q��k��X^^~=J����`�M���e�L�9���7�4�<�#G^[�Tm���y�w�K�0Ĭ!�Mԏ�C��t�:��~&����F���kN�W��,�{j�X�Bvz�=nO�^l�2O/���.��t9
�۲D>�9>�]�����hsH���%v��V�݌��-c�?h�}��h�
�B[��<�������c�AcA÷-jek��"�p=�A������64����V��|2s�A�s.�旑E��js붖nK��f��?�=Vȉ�C���)ᴸb:��J(�W�9��|Hh���4�!%�p��ʰ�B#-B*5����=�_�{qq��.{�H�����X�������/���5��%�������K�5֗��~H�խ�yl�-�3��>�a�H抃�C_O�~��ˠ��arP2A
3�V���@���&���:�K�x�����E_�_L�a�zU`�_F��+���8����k��5^�:���($�N]&����SI��� U�j�±�k��h��J!�66�Ї��M�	�8�} �O��ϟ���kg�i  0�_��n���l�˰�����k)۫̄�m��?���.�ޅ>s�a�E�M�co���**^3}B;�\�G
|~uZZZ���˛ߨ��͞�=�[��h�K*�N�qb~�����@Tᦣ���
�W�e#i�ND=��\c��GK��7�<ǚcΙzx3��'�hqY�A������Z\铓v'C\��3���9՝��%E�3��i��Z3[�#��-�;��D�&�|___,a1b�DB��\��u�~��T��d23E����9	Kn��c��%�N�n/��VU��k�Y�k��(Ґ`�%U,��)�鵅c���=��R�P �G4�;�۽�+�Y��[��~u���Ի�\;]��]��v��U%14����Ǩ�y��	b�뭭�ϖ2V�vd(�>2���.¸ۿ�J��UZ�ײ�@����C��)~��{.��g׽���sT�����UU0o�?��8�_�Z����UnQ�LNN�MǧO;&K&��/h�YWV6������E��Y��G�e�B$���zn���K���l�<o�CF�P;1�U����yK"���<�,�<Fd-E4�i� ��Y�j�� \ԏ>���ٱ��x��u{{��~��B&�{hԙJ��ȕ�ohU}� D��?t9o�Q6�rii>��r���/�qg��v�Ѝ5�������U$�b�Kf�|�(�x%���w�>66
�?��/�"�v�yϯ��de��2�е%��@���qr���$F5�1	z1[����e�]]���ʪ�����֜ԏ8�(��~� ���sysK����&SJ[�SYvv���]�x���s(�U�����?����n�Q��by�>5'�+��?aaa��9P���Z[[�R�8���V�6��CR$�_��tEKQ�S���`��e��A���s� 3���c��|@�/�QD7{�ױ�7�eL�ϯ�����E�{���`����ٙ�4��,�m�k+�}ܧƤ������dFƟ�����uy�min�SYd���4�͝��;�\�#�@9��W{�:`�zx�Wo1��վ{��Nx�M`K��0��z�uȚb��~;U�:��G����y�>�y�A�8P���ۋ�l��6Ŝ��G�� EEEe(̡��Qu��畼?ޕFu5�.Cm$f@KEb]��I��nC��/I�]���ᜉ�	��^��111`��ri �H7~�d���KY�:%������7IY��ĵ�$���9�Ž]Q
�Lz@��y��R���
��w�WDcZ�K�~kk��sR���T��(��2��WVZ�U�p�ޗ�0O�R����YJ�h@���oj���WR���YY�����)0���ͥw���S��a�sW��(�=Ĝĺ�+��:;9b���MV���瀨�)��������u�I8�I�s�֠4�ځ]����xJ��skj����0���Z�^@�o��;�"pl02x�-�gve-88gZ�f�~����/2�ɉ�\NLLLPH�Z���.6��i�M zK<-�:����s������Z����=�7R<F��A,���IO��a"CjL"��E�R)p�����#p�YB�j�}��{�h���!�G /X؈KU��vB���Av�9W�g��uujri4�����^GaH}x�&�����Ǐ�}�� ��G�C�A�xΪ���ru[U�l��'[3.�>]7\�Ǔ����u�>��������`��T������|�9	�{z��M'�N��\N�|E����%�1�'�)��f��/�Qx�tϔ`R���MĊ��w�~Lm�f�+5��CĊ�l��*�mi�S�e�I*X���r�8k}Y����p�p5��sݦ�O���M�%���|��+�}}�<���X��g�uPH�6�'�أ����g�w���y���o�Wh� �����|^�6�¡�������k�4'�$"�b�X���<������9�g�����]Z�=0�lR�^+A(%�,�]��_j�_�{�Ճ�j��~>>�h������*����AyF�ܺ�Z��u&���SQq�|�r���3$5���Y���3��n��� �������6b# ��1�G|w���� U��= دP�;��s�.�L��.��M���ʻo�(�Cg�� �T��L�yS��@�|�'�~7��`��Aon`��wȐ	@wM���ߒ0(s<Iذc$���.*ػ��Ƥ ������%�2�F��`�-	�A�~��j��3�������%u��[	H'��s�a�ڵ�f�9�,G��i����i����>�ַwpЄ2����X�a

B�댸Ujik�Ր�7p!� ���m�:?]�]
<\[k�ض[�����O���v�f�jVu�a��G��� �p[@Ʀ��aH�'�#�}H	*l��?�*�+RZ��9���-������ʱ��?o����YS�u @��z��j������A�h	:��*�[3�o7�(c\L�59��>|XV�A;���2p��2a���U�M���A�o&o<�.�pd?\��n��ek52��1B0��)��p������q�B�;�Vj�ف,��fe(P'Ooog��#��?W��ϟW�8�v�ߴ4⍃���(�|E��[���ְ N2���(>�?&a�f��Dt����Ç��zMJ��	#��oIpqsG��W���&cX�~��գĞ%�E�{
�A"zx|&��������cccP�_���]@k�1som���Vr��x㦋���kk�Nõƀ��H�f���#�`᪕!?P���%p�����8+�:�ekvv�h�Le��^�g�k��P.2�ձM���90�wΰ�"�Y"t\�Fy�w�����@�w��̴�p���h�^	�(�� :���f�&&�&������naq�X��N��/n:
.:
�5Ӟ-EZ��و���4_"�8Z��#�)����+��g��@�C�l]Z*<( �2F��e�/�{�N���q�*����7p��<m�t�D!�o54���k�wq!��YU=謭��Z $±c� �3�n���~p �M�:?�z�bY*�Mcf����rn�h	{���%j���89wv��5xh��W����y���������q��Ou�5g��!ii(��S���3��/�9�5�J#�/⣍��!�31u���>r�C��ݣ?yR�=�<��P�R���\�w) ��^(p�����2���9~���t�.Dc	^�щ!�=zgz0�8\3�v�Y��u*�����9A�}39�8�ר�Em�j�nnnNMOR��Y���mh�[U%���M[����kG��n�9hkU��`q^YI�#�%>�S�ҫ��Zr���
����g�D	�|���g�޷o�ǟ_��KKY����_�4�sRG��ۻ�����ghz9'?_�['����ܝ==Y�-��[8d���Y�?�X��Ç=㗑?����S�;~0���7��,�>����أ�:�L�2B=I*����ZO��������U��oy�2�Uɮ.�)�$��Ii��CKa��� �Ǿ����
rgsw)�"{:Y^]�s*ZL\\�9Ǐ+�І��6� ��0���G�}a�c+��˶���SSS�SCP��"`
v���ay<��!K$����fp��&JVb:ğ�B�B���Ag>)L�w���� �������'/�xH�4��Y(��便Bl�TK`�h��:��*��X�i�|FF3p�������q�|����*-��b�J��|} 'Q��號bd<�o��ȷ����]����;Q������i�!&h/:��Ǭ�J��ݞ&���:�Os��f�?!!��DDr�I0X7�$B<c���n鹼��%E��Q�AL�2��*�S��zϗ#�����:B�7��>Wɤ?u�s�U�e�7�����F��o�^^^^��yS�=}��ȋ��xZ������� ق��*I��yH`.=B���'�,�r���D{����ث��Ej|KK6}����Ȏ"몠X����0U�$ǌ��޶7��+�"&ְ<'#����K�������Ի�C����)�*t�D �h���9PM�ܪ3�va(���f*݃��7E���t�Vx6<��������;���j'�;�p8�m����ϐ�JSGL�򅱒t��U��NN1���4Kl�q����$I?HUnG$�Jؚ�x@�e��^�`��u��=`,�7�\��6?[��!�E������{���t��4`X ���!�<�NS�~uV��+��W��d��Q�̭�P��/����� kD�%?��ohٶ%k��F�$��kf������ཽ�s�TWn�E�A!!��o7��yf	��Ş�k���v��҄��3~>�Ga�,�DaD�U2q�j�b>���Ô�\��<�Natx�J�k�"�]]]�..��o�����":���~t��ڒHJ\!?91��*9tgUV�ࡀ�FE9��(����(���5��������H4`G�`�����C�[�h���X���a:EV��ϭ�-0��{����'��v�:�H��hiI�pcHJ��Ȗ�N.��Y�����Mԏ�O�q�n)*�_u���9��� ��0:�IM̌�#��F�����L�jռ�G�s��aSH����4�ݍi���@���o�.L=�����^ r4�����έ8,Ouӎj h�g��߿�]�a���rre)G{;;u&y�g�7�=��|
�n�ۛ�h��''�����V+I����?[�����$����Yp���Х&}q��;F�y* I0ߏ���d���Ǵw�.��c=�A����E��[�q=]CM�1K�A�߰����ʃ���Н׾�<]�:*�����a���J �	��'����y������9<(��FJ�6wK�����F?��]�S�-� �7X� 3F!�i��L�ݹt	#��w�''=PU����B��EK++�puH6PC�xL�km{\z�c��]/�#�]DY<3\g��gF���#���u����3?>�sEuZ����s��[[�E���Ԋ��0z�m�P��P��}��J������eX�������bԷY����,c���"Q}a	z�҈�1kB� r��M������A��� �6D Z��\�H�Uշ�04��?�ԦV�81�ʖ1of*�7S�M
t�fw.��_��)�el�mM������,�($j�	��Qƞ��ݭ��a��K��1A����kʘ�Z#�v�cd�WQ��O�"D���,
ʰ�BK(��&^m�f(�����v�c�/0v�����ۺ���g�ߑ̺�����|�7�09��]!��LPkOd�#j��D��	��A�*�/�9L�ǙX���A��/�3��)':�"g53�KKˏ-��F*�d����Ff��ؚkT�&��ֻh�D>��7����>��8���ȣ5[k�hyճ���6E� ��>�6(��ԑ犿�e��=5�3�9�����f���X�]IA���C0����_�@�A\����e-z	����/Q��� �|$����:��+W�i\ �uMok��k&E�=�7Q��ϋ5���`��i����~.��&��f�w����>�\E�Oz�z;�.�e&��V�j����oq��G5ѰWkz�cx��|v.�>��H��[�2O�ݽXk`-�*�� �֝�Nr1��!�'��?7(s�Gqk\��Is��CL{�1�x�a�Z���ZP�a�w�/���h�q��m��}qt���e�������j�`�p���+J�fDVm����p�n�	(�0�����ç��.b,ht.����7UPb��[�{Ṣ��䄺@�N}�-EJ������`�h�6�K�v�DV~~7��[�	@�ܤ !�+x���]�w���u�&K��@����ۅ��ۻ��8�r�@_��b�ȇ�	�i��nG(_mV�p@�߃��8���C��]Bc֔��%p��E�H��t%�_�e�AO��o�{N��P1�E/6iq�ߒȇ"�*��g��7&slQ}��R�#�� �E<�GHJ*�-�G�W�R��^G(?�C5~]CC_��1������+o.��u��6��ǀ�K{�����41�����:K$�X��M�� ����t������5&��d D�)��CA�P�����Ѧ1��8W����i�hU���ap�-�������|��]�or삂���W���v@��ywJ2�|�W�, �6����l������C�@h����c�n�����}���@��j�,����N'�)���{����Ԗ�Vj��
��<t$�Y��_��x������B���H@h���MQ����~���!�;��O�m���%��<_X�9�"�!F�zD?6��u4��S`�$F��F���(�fc����4�d�����h+�P�'EQ >���#�� ��A�P?�I��eU c�{.�.����#������B�^kq鴙��V�JKK[[.�B����S�l_3w{�1�ԉ�J!�P�t{�v_���0`ǨW=x{ep�1z�y�T������n?�����&h[�pXt] �h�I�$S�pKKK)<(['�{kO���/�)굹�-���";���d���2�~��~(#�3 �zP'�	h7�\\ 9�����ugT� >��Y̨�3��`҆lz��*2{
F�dU�ߛ��	�.���l�u��r��b��
@#��
����D�)����\k�H
��MF����u}hEjf�&�v�[�A�� ����E���0�=/'G�y��|��P�秈F���+M��s����ǏOe>��g�F{�� �e�F��(1��B-�|�\��!������!MU9��{{����������l�\7�|�+gaD�2ꐉT
�¥li'�<�2�6*�e	�-1��F�7N�ҁ ��qvg.B��J�aI�a%ǼX�1x;�m�7MF	�X$&ϝ;0-��6}p���!��X�q�-c�]/�؛���53��w�Y�T�h��s�\����U]@�:+���j�T�<�QM���9�����
��)m�j� ?�z�w	qR/�&��^���,��_�T��S�4�
�F!( ��6�9� �ޠ�@?��|2���P}��J$, �;/,�uV5��\�0�?qҭr�7�l�Rs�Jhf���n.U,���)����Iw������*M��������+uۛUc��
�����#�����_��Ä��Q����~���7*��p��%��7M��b���^�rJ..����H�������(�"�����ꘑ,-� p�U�f+�i2(WUs�����1f_��yxyM��&��Nr`:A$-��4j��a�Kp#�Z� n|e%p� x��8�{�s9jm*�s�!���7���y�H�q��HzUj��`�az�+�C���ZÄT6f�Ez�,��|�ׯfb1��.
C##/���@<�x�`Y�#µ$�$�_adc����ը�ӧ����j��lS�t�V��#�}46��ꦁ���3����(��E4���glчQ��%��IU!4mE�cS�[b�B;������%)�$wb���m.dT練IU�F��4�C�;Qxٞ��lm�(d���+��W,٣8�3�V-c�d@NqVT�^I��=��+F�x�|XlH�|�T�m���Kx���1��?�.xr��]@�*�$ IV{�r�3:�k�ϸ�~7�\5`!�_ -�z`����������S�&���O�F���+���c?wa\�m3!R�/����
jH6�ps�oxbD̀|��UUU��fz(F"#n��r/�N��!Cfac��>+����L�aG���/��U�a���Ч17r���(� �s�ږ?6h%���1)�?�1�U�WG)	+��+�����G�2��2q�[����m��
�1�q췿KQ�Ԍ#�s��~�� :� I�=�7���Y��2�7�.�9����d��p�7R��М�F��y��@�o\"�r7&�쓤��e9
���}������P�Wi��%����4�f�b;Hߵ	y�3� �Fh��GtF,����W�(v0��޹|:�z�}������188853��C�	!3��I��9@�y��;��IG�ST���[�����`%y�/Z,hZ��NM� ��~ q�s�u=�+�l��5 ?�9iiW���#hB���?tvuM���VQ��,<,<|jidBW�^�+�k���x%�*���Eg�3yB��9�]V��:+���䐆P�(L�ʻ�����ZTPD�i�fl����O��h\�pL ����{��ҁ�{�o�����e�Y;�3��L!�G���&_2�燆T�ˬ�`oN^jΡ�T��x��"�E��Ў�D@;��^���^�RK�TMD��àD��1o\		�b��ξ���h;���r^�Z	�D�A���I�L|}�
!nA���\��!ڛ�����[4��W� �K����A�L�n����m��<,]]]�#w�;;:,�1�@k�x��F��~�nD�Х�߷$�T�B��<ף��0@��k�g�*��+���M83��XF� �e#޸�w����JlZ靆�Zs�h<۹�Ś�R��HIؚ�(�5aɼ���%cE���!�U�%Y��h�{�p)[��B@ݰ�7�����jHH�S�B�c�%�4Hj��LN��Tf�7Œ���(=>�]b�c���zF�ӈ�E�3�Ä{*ʈ2t�-������H�4�z���Z�.W���ʰ�-Jo����&3�U�}�����%(�ă-�"��i�*́�\0�T����=EO_����8mF+&&��Ƽy-�|��.דQ�>tB�s"p����@4� �� ��c}�|zk}.��7~�r��VRQ��X]�����<h��Rmcn	���KK�K�*�1-c?7{0�*D�x�ҥ����]K�H��@7�@H$�/\G�	�ߛ������堼�?[@
?;$�Kz'�I�bCĪ���_�ҹ		����?@�9��q�D�B��Zً^bI��C��Z�����D�:NNX����y���0/fg���Q�����<��$2K6�y�Ə���N�����<~�?ʼ]���:A��mCx�|C(�S�/˙2�V	E��:�ќ�Z�L'@P:�u���)(�k���x� ��cn��!��&�UU����׫�S�R�/�{����'�k�Y� I�֙)ņ(0a8A�JH���a**#�ZY����$J���IEa�"Zx��XE[;���k� � �*���}3GV]����<�1��04[1J)�Oef��,*���EzffD�~jCb
�kN��/����u��� 4A&=|M"�!reW��59�a�:��hE[�3q�f�Yp��Q����������^SU�i���
m��b�DY	�2��8裷1h�֮�������H}���gO0�*�ٳ�PSR�;:���̱}��}��� ��`�;�\ �����wq��/ ,��^WW6PA-�,��O׉�R	;%�iv�
�4ik2a�<��k_x�I���EX�z���:z���+�ߒ��Ё��F�C�m�3jM7>uz�|������������|*�!�=0Ѩ�b�NOF�Fx�)�ٖs��[?T�U� x��Mc�/g\�'!�WOq鶕Z<�ScBL��
��vu4i��u��1�:Z��#�n]�e.��QҠs\��Sªe�0����G9`�3^đ�:���e;����%�To��c%�2�QR(�Ch�"�<��)�H�2��IHu��d�L�#!eH�B2d.Q���C��߿ǽO�:gkx׻�^{o��n~>��d ʮ��u�� �&�����`0����u6__�=B1�>��2\k����v�����p�@D:Gj�oŮ�گ��|(2�2��7߾=����'�"�e�A�I�K��@�Y�����`�qf�YY�Cʱ��i\~��&�_1o��Q�t������\��_����{䨪�<�QDx���ȿNnT ±L����6��?ξ��k�(:��^�j�Z�Z��H�~�9	�����9�~O $���}���š|7X��Fz����>'�yc�b>�)[�����]w����pt~�/��?�E��|��n]�n~QӏO&
�(w�C0<,Xq������\�"tk^9Gc��e]��{��B�/1�va���x�oh;�7L���ϯ�a�{qm=�3�Pm��`g�|� �2�8:�y��O��1��E�8�2���_s.����1�\ �~{�{������WRi-��;�O�� �*=,C/Ni;��j�y'��߽Gߜ�T�4X�� ����\��~����?ο�~~T�oq�o Xஞ?Z������l�-�]��Mk���6\�Yl���-�/`��¡��v"��z/�+���1^�u�!�r��	��3��(Zs��,�0�rL�=��-�j{��u6��y6Pd���f����$�g�C��J��>�+~�C~zE�i�w?�~��º�#G9o
(m	:�2=��ȥ��3����Ą��rS8��Eb�R�6��M/�_�_��і�Q���x�Q@�qq*+W��vÎ�1n�;#w�Uε���������r�^j��a�!�5��=З�dR�ҥQ��ĝ`��A
(���� ��I֊�.n�ԋt+r����[�XPH��+w� @��#~oU9�	���4���r=<,,�I�p����M��׿[_w��n�=�z��b��#u��#�m�_��f+/�	{.���ayG`mO�����&�e���U�M]����GTT0(m2���jd�H�,m=�R8��0�� ��|�9/�r�i��v��{��&#���a�^����c��=Ƶ�cƖ�%Me�l ��!�3e��5��SЊ���T�Q�\ �����Q��!��bCu��̻��¹�/l�����:���he2�2�x�7+�GQ,�����\��|ZȔ���_`���7���9�+�:r����ߖ�"�]����Q�yY����q##�OȽI+u�v~�6����G [�^x���X��p��-��m��{���z{<8�p��sO� ����������p����B1d, ��0�*@��ó_��f�@��4?�V�qz%IU͍���j�`oi94 &���D����RG��|1�X��.*�@/a1�m�D���eהk�$覴)����b^)[/�:���n��(�������#���
�Pz�Gutt4��6t��?���yS��&��2F���� ���ϟ?ҹI2��U���C*1�&?�/?��B_-n}t�-y9�,N+m���:Y��Zt�`��&x_Z�������P�U><\)���*������9B6<i���^XT��It�M�����`��G�_��{������s�]ʡ`��X�ƃ�ې��~6�6U���������v�����|b�tXm���h�6Mk뎴7i�e�1�_'s���������
�>^v!ݼ�av�!D�
H&�:?S��Ӄ4�OB�K��z�'H��]{����fF��+�Ph�z_�C�d]n2A�__��W�j{�h��8�"��r�o�����}A��3��Q��m�6l��7 �p�/��'�]�g�a�em���n���Y��{l��yI�0o�}��̸��&���o�kd�U�`����E�wYVF��b�g���싘��j�*߾�1�KdR�D0���e�_����:t��r*_��Ҽt���ކ,��o743���Դ�W����P��@���W��� L<��G�.�&'���	"�p(�?J0���@t�	d,�?��+Cr"|�a$�BƤ�8��ɚ�ˆ���p�ݗw��Y4jjk?{�����i�v��ޟ�x7y<�,�E�m�Y�O�6,�/y#˕=�Z���n�|�BB����.����ĉ�0Pp�-`6�:KB��7:�~<��ڟjQ������"}!�ئ�7T�5Y"���
	�M9�M扺 ^լaa�T��o8��M/،T��w���놆2�y'䖵��c&�,N&^��-W��M��*�q�+m|l`�u�ǏG�u��J066�����%d<��2;����nA�ϐ��ٔ�LF��#�ƪ�� ;��@,ܻ3�
��5x��K�`*�m�����4���32R�&|� W�t���܄D�6�g		���Y��#�4#�:]����lxvGv�����*��Pů�eN]j��/�~B�u(�����9�D�l6�khkG��jI[��x�L��f`]7�I.�����p~o�������6-��X>k�Һz/�8�YE�ӧ��c��4�͔2�<��]���ǚ�����~L4J��
�r�Hw�H���X[��q���T<�ܐ�Pfr|���(���{#cno�s��;&�n�wr�������*�z����N�AѵL;_�8�������Fr&o��Vsf�ǥ��_��ʲ��Ns���*�Bׅ�~]�/�tL�������d։���B�v�7AWrr�w�z�GeUՓ���@�jsv��p������l�H.�9j�j��t�=`����A�w �p�T�u��H6����p|����^z?���O�t�k_�Z*�:9��ɉ��5ww��9�ZL1�J;�
2�����艺o��z(��'_^� �p�4x�*������s~w��F�P��!�d:��G�M�����¯�]w�J��B01�����"1��&$�z�����6(�Ι~�S˛x4�(�������79�̴o��Pr�
��g�{�%�M��rĐ k/E�{�#\ggh�j�g�iQ7.��5��kn缩'@�|llL��`����"�@G�ɜW�Ź2���E&�MK�M��?��:�����A}�'~�;�I`��R������h;��{R���888t�?����^���ɱ�ɾ`�9jjiu���E,�������x|����rSM��Ǜ��k���e'K�P�L��y.�0^�U,P���j�U�����ɜ�Ef�N�v8+���n�[L��)+���p}�js�l�R�����C7zHQUՏS��)�����+B2�i��T$�� �=��UP���*��+
j-�Jz�v)�wl�������b��>�X��׮��ݵt�>�w}�a�9�5�)�1�eÆ}��K+ǆn�q���2��[2�&�#VC|۳�=t�Л���A����2j�j���6ۏ���]#�c�0)V�2|���Fp֔����,?'��ԏ����1ժ�~E5��Ɇ	��?�	4�2����}�`��T�|}}G��'�����(�'{!y���F��Z�j�,X O�O _��Eb���	Vk�D��8َ����1R���bd��e��w�T�ģ`XR������g�T�P�}$fQ��nk�@���j������h�		5�j��#���/�p���M<����Yk�yv��%R�n%�g���U���ޑ�����)��(���2|��]�T���T��ѭ��Ј��\B6䓊t�#1����[9!�c�&Mf���ڴ�IN��-<���t��󜤶J�l�xSW��u��k:t���V��F�K�n#1��߾}���s��#p��t��X�_��ű�~��:K��&.�S[�G�jq	���� p��T�v<������G]��k�l1�63��U�d��6^J�)&��b�הzQ?x�#���ֵ	Z {������3�f���D	II�H.J�K�5�?��*a^L=��!oN#7k	���M �p��,xeޒ�/N_�$�G3���iڴ����WQcc.n����������}�f���@��ޗ�'���{�]@��A��=���˛uɚ8�N�������K��`��|�B?�X,a�׸qe�-}��*��j�����)�	snY ����=�s���W�+�5c�P>4��[ׯ�r�W[]�{�#ŚF�����V,�8�[D*X��9H���ɡ�U�l�:�>���������������g��}ddd������
P���-x'�=	�`�CG���cV#������ݧA�:^ �e��`��K��5d�		)ӯ3<p�S�����g��;LZ��� Y]m6g�w�y��%���nZ�p�YCPx��� �����"��=�@&TƦ��G�eFD�{�y���Zy#���1��n4���=��Ku��F~�OƝ�9W�w��~qJ3-Z�î����/پ|�Y��	�Dq�����[�frVX��5��C�y��O���]����n_��v��]]]5<
&J��B^:���u��Z��$�L���|���{2N	�rh��ƲiP�R|a�"�����@ ��V�]��ȹ��R7:�?�a���ۛd}g|tT	�5��ԏՃ��ѵ�U����V$�g��`���4�
* V�y��3o������q�_B��whA�'<n��Ө��v��K&��#�*H,\M^��F���;{�g�$k��>\
�s㤢5�ߊ�5�{m����>��>�N�Ie9'��&��U)��E���#����3T��o��]Z��o�G��nDMH$.�9�?��i��2��\�p�H� ��y�y�*ס��5<�0�������1.��ц�@D�]�+�����6�����h��x>�F����O@Nl�Ui�4-X��3�^^�]�^GXL:�u���X)�4ɕ4��/|O)�O*H!���k�b��[#=��[H�}����emR~s���N�R���#���='w�.�'��4�w��D�����]"�����"y4>r(�k�����$��E\�		g�j���Y
������B����_��𥿽ie�WXX��yi=jB���Q�@����V	��9�� �l���0������'%���x��#��> ٳ�b�aӏ������u����8�<S-+��j������ey,�y|�k�f�!���\BB���`m���u��c�]- �C�ŧ(/]�x�cﬅ������-JR����a�=֗��j �;���Ѫ��n8�.u��ߥ�8TF�K]]B[��'���V��.���W��z+�}b�����B[���K��ן���KKK#.iij��^Y���P�5��OS�ֳ70��c	����ۮ`ۊ���Aaa��˱����{�V�M�5<s�A�z���_����t�O�������p)��;!<� V�P�<�'^?���%k��ȑ��uN��l	��V3����g�"�H��2Ӧ�6�U��C�?�v)�;�):R{6������X`\�4#���U&���&�8��s7Y��ϒ����Սq Nv�r	UF(�"6���h��>.[|�#��R7�b 0�K�ܼ���|1Xb��$99�y'/9��/xxP�~v���7��ߗ��_�!ر��� �^GȦ�/	�8'F@�7iD��h7����c����F�%V16��D?Ö:�ɇv��}��gz h!YYY�8�xr	��'Q��A0�81
���3�q��ڼ5ܷ^@��%��[�"�(^h �8W߹zI'=��d̩�$H�0����_p�ׯ_0l�7���m"��R��X�7xpX[Z"+��l��p���q����l��H��ƾ�Cy�쀛������27��wCI6��[��b$G;t�uyrŴ���&D��`��CDt��2���DF�_���`t� ��������IwVZ�QQ��u�^��AgXH�蛬�G�D�!w�n��������	��3����}��$���M��}����%��?K�0����w�Un��ԑ�.w�0�~<��̏�4��]	ET��cX���X`cҰ��(qXY9�v��#���g�%?#��� �a �n�÷����XƷ��� ��IE�MHa7����n<$-l�dݯ���/�:���DA���=����g;���Z�u��E&[���V'�8Sm�D˭�؁�`�NuC�������)���y;i��KǛmR(�6.�Z0Ȑ!���Ԕ�\Ν1�inum1b�Н� +w@S���~�`���С�����*f�o�_ ������ݳ�Ȃ9���<u�N�"�X�����'j�l�v� � D�3+��	��+H�(���kK�k'�Q<,�OS�&67FI3FJ��9�b	�|#~�Q���AT��e�B`�׀w��g���!�PH|������L]��뎬>˳v0w���.	���C��� |��0pi�b4\5߹���(hC;�RL�$'��9i���L���L�p�DP� 2�s'HK�gnB��Í㞆,���s�G����YDs�D�v<%Vq��+@;e��G�M鄼��""�\��g�X��=WX���i/^�H	ω�Cx��c�u=�:ܲ��q���h~O��m��XOJ_) r
[8�	ȰZ���_*lNe�jR`u����v���`���k���2Q.Cd01][[��U4S�p���X�h���i�w�$��t��UR�2�yP�#�l�F�r�yv g0��Y�mZ~b��j�����>��lf����F���j�C��2`N�[BU���G��.~�������5�D�E�ߗ�{�Ҭ�GJ���?���2�P��2	��{عO�29��J��K�.���r�+>y�R�&pA��Õ�h���o޼�O��
���ڪ�7m�'�����b5<��Q�}Q##��
��M��
�� E�X	�Nr���̑���&�y $S�����3�}<��˗�%GBw���ɂ!�K�����@���������'���7
�c[ed�pKi�ȏ}�;j���aR~���HC����i�Q4b~b�G�}+q�O��_]�S)�~�Y������֡7ϴb�jj�g���Ǔ��	�V������0� +�.H��s��0��l�J��<�;6Q����%n}L���~Uy��]�Њ�֛b�)>���.�7����V��j��$�22�$&��n��H��8@Ӵ�L]�hUjr��
6ρ/?�t������&�n�5!����m�c��_�׳��v=��߿���"�)���J�5iZlx%=}W�^J!)�
2M$}�M���E�+�����&dd� �0N��|��B��ӳ��,��/��iffV�C�Mț�:��:_�ĉG�E�%͢�C�g��ӗ%fER���p�3��G��Y��%���,�?Sx�"��`�f�փ?����ſM�CDV���`���0'Q�E�cz���㫿��T�hhh��i�.�K*���}M[������o;%����m��pVٸ���Q:70�¼Yl1����� ���g��c V�x��<o̴���i[��2B��C���Ϗz�V�$��OF��e�3�9w<	YS�=�2U����|�lJ=�y*�71�1~��72:��sr������ѩ�1t;��#s>���]�87���oV  w�!�+���(�f���Z�RF9xuﺶ�l^ o<p�ӑ�I`EK�qi��.7�,>E
��I�F!VB��{[��֋vE��d����5��x؁7:�.�x�0P7�Q��˗x�8�Ltٴ]���F�Oj�)E^�/�9׬Y�I���	�_���G���2���`R>~��~���y9��MC�3g���l6/�_�b��mp�	-#��}����OX�RQq�zb���?@��C�-P��4��:������iȬ ����M�r�[��b�-�F>4�%�@��&�v1�犾����Z>*������~�� X��=���)7�v���������n��o+�ș�^�Z_oM=qW���ǉ5�H�Uyt�-�IA�>�>B__�G}LK:5�̹M�! tOO_��ˌ=��eۻ����Eݥ
@��<��5�u��ub-�T	�B����x�=55<&
#�Rd1���
�i��JBN��0`[�͢^J.$]������(xCn��9�:̇�+D>i�ֵ�T)��y�Y{i:�y����ԅA/�V���I�K���d3�]}xs���C)�ׯ�|�soI�o }���� sC�+;�N�B�OO�� #������[@�h4��:����dރ�: }w�|�se �e��zhL���!���X�t�ҥm�� ��Ӭ���jj�D�����\^��Y~���L���Ԁ�H�8��ׄ�6 o�$i��Ջ��q�s����$9N6O���Ҷ�������������<����wG��ځ�� X޽6Z���Gÿ�|!�f�q���]Gbb�y��GU�4���Ŧȏ��wT|���~��� d��D�5A\�g��V�gu�����6��>%%%�E;33�Eܐ��?c��H{j�,�"c��ͧ��{鿅?�,>^KO/��4 ���S�!��].$��}&�KAwvԙF)ρ�K���Z<i��;�k��"4�����Aj9��X���k��sg��[�f�e=�O�EI�x��9#�x��F��۹��S���OLO�nkk��g�/���<�o`�D����Yk`�*⫴pה��~�Xё���ӬC�/�,;u/�� �gΗ������ƅ���%�&��a܄��@��w΁ �޽;\]S3&��x��A������MP+�o���:}�	 ��74�Lc��Ç�{a�sO�����i�����=��-W��t�}�(��!�ce%�37���\�WcX)�/��;26%-�4 >>P �T�rz�������x�!l�����Ss�˚��M_� �Ά0���Ξ?}� ��,6��i���U���NH���(�Wd�n��� �&iZh[��*�V�Ķ��ŋL��hoN�)	&#�2�k'Տ�7-���3K=>&���Ke��v��%�	�K:�[�bKEm�R���M���n�o�=����?>9�J��$�my�������iI�A������}e��
S��R�E�w�� �u����G}F9i�����"F6T��rhh(���wIH�� ����R��b�r�.�>S|��`�%�R(����݃37 �m[P	�ھ}W�'�z����P|{���F�OD�G ِ��HL�E�����p��8�$����Iv�)�3��H�,OǤ2����pIl����"a����C��N`\Dث�}}*`�M����;��׀�������������Íۍ����(I�!.G��hL	�`�QDI�m{G�Z$ԗ����9�ӴӦ>�����a�_k��R�@h`鎌��T�@�"0�������+^�)�潸Q�ބ!<OK_��d�]�O�N/y�h��O�t�O���ˊ}�K���q�΂��,"���=5#��k��U-���N���*GV~/���?s'sM�`ֱ��^���\�깐�׹�x50.�0Q~�3#�&���v�`:h7D@��Ǐ�.Z�$ X�0?�Y6���54.�i���V�^=gI�� �?}��|�x��*�w$&)y����=���###�E���v��<�v��6_E[����P�?AF�ٲ�a ���S��=HMo��E����]�B`A��f��u��=z��s�mii۟�F��T	<��1|���8;�XT�����HC���f�wgg�z�H��7,S�O?�^&�4�ge{�����/y�s��u��i�sg��^�L�#0�C#}�K �c�R~��e�"#�*����[��k�瀯!�R�A��Α�D`¨`C�7/�SE�|��W��(�����{&��<r���R9'}�����2-6�u�2�>\l�K���b#sY�� f�VF#^=o'�'H'�*�9��n�Ց���a�Ϸ?c�O�q��*�#S�������^F}���#h׺����K�g�P&CO�0�:r>�ii1qq%�Zb�����kJ3;uʲЇ|y% pPv<j:��
�f��m�ٗW�#X�a������ů��1m�SX��9̲9�Ep��*�]�:��<�Q'W��=7�pd$���;�DcHKK�	 VU|��sC�,�4T��Ĕy���P�X���f�Lu!���)y!��S��l���O��� �F� �� 	�Ωz8�����Ga��(
H��)��ɉ��4����E��T�Y�p���M�=�஌S�@k�v�'��̮�*�z����\�I�V��{a^��*�j�@qկ�<��U��<7��R��:	��%ȹf�Y����O�JH;p,���[G��r/t�?�Ek�|I	��S��ZSw4��'�{ׁg=��?��J����C��ҀSXO+�k��w��ie������0�u�%����OwW��$�2n�U与�Y�cl��KVU�­�}�����ѪT|�������E�����P�*X�dA�^�禔377ϖ�fX�>�~�L< T	*�!s��VP>.���jJ(��D�h*$ `ٍIj_���3�]��^YWW7w|'��v�B�)͗OF;������t kb�wn 1(-о��j|�����7�ֺ<��F�<�*�dFe2�GC蔊n���o\�(|z���0��L����I��wt�Da(���K���zD�~gC<�e���t�eй��C)%ϔkr;�e��`ֆ�'��O�fFm&E}��/�hg�p���[�<��,�����/$��0�xb����}9g𔨇�b��&�X�kC�r���n}S�ԿDLtai������kj����������RƘ��3�����9���P�}~���uS9Ӝ����h-c�(ط������
d>~���`�u^�6m:}�L�*�Ģ�;��3�����x�᠟��T�=>D_&�����jp�,0b�����ɏW��H$�&�<�/�j�6H?Hes|
qP�eͬsQ<4��9�R��K��;�j�#�����',��ڦO���(�ǎ��6]�k}
����]YYM�U���?6A��р�I��<
�]Fb�,���y�hO�q'����'/n���75����.�b��J�HB�a��8�}ۄFA����w�ϟ���N���9� v�]�1\�X��q�d���o{���|OO�±��S6? XM{��(U�3Ȁzěn÷�|Z� \Tf_��Aa��~��Ã`��Cŧ~���ߓv�2/��K��)�L�{��,!s��Y$�S�	j�1Ϟ�c��5��ꘄ�Ւ�Uߊ% �D�b�H�"}��#��A������� _�w���`ݾ�+�WlV9
#g[�0����O����ir��������s��s�!��0���yE����-C�8 Rn:,:S�
:���ӧO��|�x�1�}Hc�1�.վ �A!!�SChӁ�1��l�`o`0���RWD�ْ�>_,|a�q�=6�,&������D}N�(-qѵtk�|wA�����b��H\���Ш�u�m6��pnb��}�Ԥife�ڽ��G�z��-��t��b���ׯ��Ret$�#0�\�8�1I��z��PaZ�=̡Fό����x�YP@�	*�Z�{���P��|���|�w�ڋ����;�^rs�1/{*fq��u5V�
/b&#�c�=D�>&��2 4��(]p~�+Ȋ���K*k!X�,���A_a#B���޽{��ٽi�o,�Z!�y P�.lV�����d��ƅ����ץK/!��kP�4��-������E{v��$ǭ���t���h��\|��5~v�E�Ԟwj�K��K�����Y�VKHa�
kc�����C��P�/�����s��B�I��M��ÿt�ط*	��s�(���2NY���|r.wg��&Ar���s�IJ:�{���l�z���F�/4��<�y7s���ظ�S�>���TFc���? կ�B+Q
PzCZ$XN+p���_MuZ��`^FNN��Q��b�'��Y�yY��C��\��N�)���>�ym������;�T"ы�K�s��5�5��tp�D�/�X���N�\U���� ��a��@�ކ��[�</�\Tpr�Ԣ٫�F�%)�r" @�&ا@��s��=MMՄ�A�=v�׊���������}�����k�)�i�O�7|rjgq�k��@��R��&oo�̆:�˄�T�7����ƀ��c����]6w��-y���D��=x1|um��P��ġ��xf���	y���3u!���߂�0�z��ΰ��|J�w��4�'�ݕ� ��	��Ί��~2s��lć��
`��ҀI���<�|�_����&���\�|�1�K���)_�hx[��Y�V�*J���>��@��z�Cw[=�F����L��xtߑQ�����߿K s+��c߾��T�(���	n�~d�6��qL̡��x� �p��'�)���+_ZZ�UP��`_�(�$�Ű4��;\��2fyio�}�I	�������c��s�%�>�i޳kh�df�dfEu.8f���57�]G΁���U�1w����y�y�l<S76N,+S�a7ܜ�|h+�9=��x�O�8 FX �
�L��V�b<r�'q��)���>��^�"���� ��8���C'���O�뾸L+���QMh�����'��Sċ9�c1�l /�~����LPLLO@�W�]f�I���t��˗+���r�M3��=Q1l��:l;���` �X�2�A���3�#6��a��T�Wޫए�K�����;��-�o��� Г���p	<s(	UG�=�Ԣ�lܴ|A��u`����Kxf�ˬn)m��'�}��O/ߺm����k\�(�8��14�0`oh^����'��i
�>���z��B���w�p�pN�v�� �m<�>}���ns���#)�X�︊���=W�E�B�qW�Cc���L���N��;��|����lD�ٖ7X{g�	�IO�!1V56&�?��O�1�}������N�$]��r����:2~�������3�z%D?�B^'7:Y�k���� ��'b<��l��S�U#��q����@������EC��!#��C��'ΑU�*��ij�k�4�i=�8���bA��tڿJ�KZ��� ���MSȾ��9�H�RL�b	|����/���ȿf�^zo��]j[_�H�j����½]�q���N�'�2}�i6��c �rǁo�+)IU�׺Qp��3M_�k�y���̰�:v,���M-]ݧ�M�:�[�7:Q��!1�ͽ3� �½vVç�I����G%�����p���_�P>22R&��?��P|�)B82!���df�g�ͧ�Ok�%�~S�����)�|�����f�����>&�|Y[r�������C^������43sjǘm#���ϙƾ��OS��%9
 �⫪c4�����dUWV�_9�'���H�#�e���0':����y=��@IԦ+w���#�Ꜹ�FΛ;�����.~����� �VS]I���W�;S���591zo��7��J,���qjl��*E��9Q3ā�z�P�W��c��pU�L�x�=	嬬��!.$���X`V�����O�� u��)�z�\�#��E�@�1�GkZ�[tlG�, �<Р�M������]��ծ��Ճ�^���4��u�j%��
�z*sC�'����)=|c�!�]�~��%B��|�Y�zW��ĝq��p��[b}���EZ��˵����Wd���*c=cUF��w]�Lg��>~���<���MWel:	�`��S�l���`Π;w,���=q�)a� ������@X(7��#`�a��z����{��5�������t�]߯���+�q�c9�oii���,!1��7�
ֆϝ � ��RO Bifn�=l��x�ڢ�Qh'����6l��̭Ӛ=��G?�
�C
�s�����	Z�l|�������l�j�'0��K�cuM����;�Ұ��_iS4�cJ[��ǋhZ  j�U��d������M�0[q��TEO/75����XS�4��.R�gJ(DOo��������5��I��TjF4 l�ܹ�[��}�����k&-~��$�����I �)0�[�Np�Fn~^��G��_�~[X��\Fo�'y���{ϥ�T���թ���=�\֝��X�u���L��c��/k8Ԙo�$�tܽƉ��7k���ڞѬ�o�! ^�u������V�Q=��*�$����<<^999o��9��HAf);�����ʰ�&�3;pz���6ױ�"��x�.[f�ݯ��?0|l#�y��Ή1
!	��5]qn�iI�5�	��wc:��܆r�������D
��4,hd�5��%s�����l�5k�=z���Pw�	�ԛ�<Pq�5PM��Qs~8��H���&G��k=�V~��%k���Z�*jk�"""pN[8�b*��	��,/��t�p��Ȟ����p�5�uRΑ�$��� �1+L���(��}���W��i���;w.�40&%�R������V���/�x��T-��z4��}��W�h�`l�SO�Q�[j��}r���(GE�%K����⒒ѪBBk݆N�ʹH���AdR� �M�T�x2lm"�C�3�}b�yb�#�ի݊b��10"ҏl>y7ٜ��E��H,O�����~u�Z�5�<��,i)����5x�'�%������/��F«tAL�I��
.y`���-xuC�9����c���'��I�^�Y������z����w��?�c��,`�.�'�3t2{����Qk���p]� <5*㷆�?sVC$�w�^�����8��|����97{vvw{WTT覝�*�'!�XWKT4�L��eR7,=��/�X�f�*�	g��o�Y�8��r���-^-_'~|��tU�����h``��qWM���Fe*!�[*���}$�}j������|���S�gL���;�:B�DqH�_������Bϟ;�������Ñ�ݩ�X�/��_;q4%
S��̛���*���e�r�6���S*��Wnذ;|�������mt�Q%�$�f������[K�^������jM�8؍eY����	���sr�'��=�ÿ$;@%�!���]�}���t��v�n�H	�ft�-��ڧre�{d�Ђ7d(O�(V��Ek��c��ݴ·0�����7���@��������,��P���ɹ= �P�m��[���ÿڎih��.�;;6�!��8oi��tDޕ���]�%G��@؍��<�����*��o�!F�kǚ�����8l�OD���7tfzWӓ��&1w⢸�D��G}||�<�v���&��?9�CNN.�x^���������ud/x��r��&���N��:��t��.j;/��!s��IU8+feY)�-1�a�xkME}�j��Qѥ�{O�˭�wk���+g�\��O�t['�]����F���J���h�0���?_�U�] _
a�lr������v���G]Z���/�ǃt����m��&ɐ�����͠Q�
rs��<�P<]L���U��}h�|F��P
�+Dn�/�j�-�"?��(�����vq"w�;Rޱ�"����'Ё�}�~�Fy�OmY(��j��lrc����������I�u;��
�	G�
��FIػ�߾��V+Ry�!�j@=5=�]���]�V��<�!��D��HEc-K�m,s�0��fů�i��8�
&��߉��:���������ٺ�Ŵ��-�E���ƙ������W��d�+���8�_4m���<Ϙ�N�M�s����':��V�7��xr����C?�����y/8�o������Ԣ����@�bd'0�M���w�ΰ/^\���[�F�1tL{`�<	�C�-�`�R�'s~�#�������g��Ƿ�>79�[�;�>�Ym�R��%rw�[�~�N2R_�T�E���g�5���|IFfr L����^J�p�tG<����|�3�9:�}���u��Z���u�GF�ۀ�D/��| ��z�*��8�������|��h�&�D#�I��6���f�)��I���</�.�lE(-Zsi�v�!���iEc���{���@���� ���_o��^�y���+�d����r�W'ˆ�Z�[�b4b�� e�ޏWz9���HL���9�}Yפ{Wk�ހ"�Ы_oI�#����d�N��)��#$_[�Z�U?��i��1��,������ϯR��?���C-̟.m���%����x��s�T#fy4����kݸ���ϡ��bA����ɿ��&���֎T�C�n`�x�LQ�|= iM�?����/}n� �* �,������osfR�qп�5��Sq�I�GFG[�B�U�,K��q��	��L���L�Rt�<��0��.���J�po�QX�R}m��,D��L97��Q���|v�?6d2J� ��X=�r���d��5�t4��3�V�!h��X�SP�a!6���6�"Lf\B�.���n� ]|cq���o5���0
�iu����?�����A��<ΒK�½��	���\��+3!u�7����^0�-����s��A���߸��K��<�MYD=��@9�ļ>dz�3J�G�풓#1l.X~�p�p�~+�O�nW7�V���iI�2�	����$1+�WO���:3���-ɉ��ʐ�Ŭ (;[f$ɰ�gӯ¯�gct��5�t�̙�`Bc%�S��%��IXkc�>R��wf ��i�Mˣ���	��3-������6�d#��m�xӔ8�e���;,8�fz�.
�м2��9Mgr�^��n{�Gm�����?#k>�O�:X�ŻThsٌ�44-&TN5���?��孃@~pG��.���NL�����1�Y�qM~�m!��٘�ɷ�'��j���8�r:�X��N��-�m�8�6$te��*8�c��FAo�m����� ��0�6�XAw �?�?��؉���&�R�=�>h�cin�8	���>TU������9��C�2JvLq�t�m�BB��?���.���.�E�S������G�SI�0�L��o�1�?ZH엚^~P
�<���@�UZj*�@h�~��S�J.f"�^��Mw��N��5�����޸v�Z�?��@�o�8�5�8]�
@�N��2m.�Q�G��ZM�*�9%A��\ܐ�}d�1k���3�Xڡ�>(�R8[���%�	�u����V���:{�0�>�i~��a�;͙���������刍߶MM��@>�5H݂ �.t�"�����GsY �p�C.Ғ��t�^�M<�-�^�5.)����JD�"���|��
�[��L�3�m۫�*#�N6�	{'2==��^��2ߓIwILe7������y���`Fƴ�H��2*8:p�cF���Q�u�uLBB�Lt{o��8��F�X,�<s�L���bH�+*������~�.,X���}���OH��RQ ��U�s��)%��|�4E\�oC#Qm�k�;%�!օ����7�2�K�Ȉ.��6oR�M��8���Be J��dN}�FH<U������v[<}���^VB+��K��n��=߿�`�M�
�<��8�룋�ݳ�KXe���������*�Q��8u���kl����_/!V�yoA80*z�5�ʖKz��Y�g� q�hR=�����=�{cc��NvO�.�P��D�mZ�~�z��23�a�_�P�}�_2;����|�j7�#{&?d�>aaa�1�n���i�ijr-�8���!��;χ�ڐ��`�z��0Z�2A4���wV"Ȯ&N/����jz�$�
�L��&�M���眜������{bFL+�w�}���I��ro1(x���>�`��Q}��tEC���]�`dF�$(I�7�fJ�*Fjjj0�mF�R��*���zW�&4w%N7Tlkj
Q��Y�^���u}Dq�[���g9tDMk�-udd���ɽ��Aڂ'@+�b�t�F����ψ�l������қ\"�Tl�tT,�6�|�hu6Ǐ���; �@e�_��L���0X��zw�h��<�����+���M���c���] "�q�_H�de]ݪ���(�uK�O���.H9x�!��+�ٶz�� �F�������߿�  *FFn������ G��r����͞�?���l0+k٠B��X:-S�T��"|����D�=|�s�/v.;m.4���i8Ԉ�ݦhllL�hV�0���U����*�]ӟ*Z�Hջw�>�p9�������'����ʜ���b���9=0� @xA�ϟ� 5앥��sgZ�O����Q��d�{�R�VΛa$V��W���[b%�hق��B�W��9���iS�t�t�fP0õ'�"�;��A��z("��P�THj����7-`�T�ȝ�����-�M����߮�6w����/�K��8)1?&�˯US�<���\L��.�8�笀�r��g���}o�Vx�����!u�~�����L&�s!������h[�\�rl�Գ)0T	1{| ��>�aqέ��K����D���c���V}����!�!e���`�LN�.����w�]eZM��[j_�|���� ��@��ݻ�-]j�ċ��%o􊔼�n෯W==-{n{�L������*������/o����h C�TZ	tٴHX��J!��Ȣ�(d	�BNjZ�'''�6�웓�cim����677�ئ|�ĵ��7�OFc�>�Y�����8�t�>��D��<�Yjz�N���ģ�`�[!�E�K���>x��V����������@20��@�f��6��py^n��	���^��0�ǃ+0:\��o,\��ld�������t��.2�,-J"�#1�_��Ѳ���B�Y�ظ!zC�Y�B&���i��u�G%�\bH ?I.ÿp�̫%m��O}rA�qn�q��dkkH���00�6K:��_XЊ\~��[����n�;@Б`������o@+��s��n�A���&e�/����V��#���zմ���@}l'��K2ՀM��T�]h���O�N���d�v�a�" 
>�� <�M��]]^���0��ջl>5q.�r��-��-"B�q7����P#`����]�adOOߗ�S�&4�X�D?�����|M����>}�E�_FP��B�l8<�s���u ;��e�>q[�&����x�A=��"��í��o��ˡ�r�\Ļ|�s�mK���F0P�B��������bw�������mWˮ��7f?D�gF`X��*`��l�Rg���:x�D!�� nr��6�7�[�~���g����-y<�a3[0��n��>���Ba'k��e 	�.��\	����I c8���L��<g�i�b���zj2��́���2A�b�o��6NhR�޵?FDX̝��4-��)�MgO�?o�Ic���7���_��Jy����jժ�66��R�2N���v9�PyT"a.��k����\�����&�
�B�T2;�S���I�<ώS�Dʔ��$���n��3�e��3�w���������/g��s�^�Z�u?���¸�vsV��0]�jK�=�qp�p!�9�����\��$r����� ( a�{Q^��"�9J`Zg�WM1�UeeM
v��ia�Imu�A�� `�/
�X̢-�*�C9R2�>�2ӚW�-��r`3sss8��o�'���]B4Cv�^^�d
8~��OY�cT�)���y/� ����h��oݷ�>y�d/Á����J��-��X���MB�~�ԃ!����u�Rʏ�J[�d��OP����)���6�*�i:���|^�Ao�|�c�Y���ӎW�<�ry�-e�Hi	�ŔNH*6t��;���A I��>\�'��Lu�&�@^���-�����wu�u�I�a#W@-��34�wY�ms-.�6�nhbT�jaT!w�3�1�,IZJǡG��:�Z�v�a�Q��k;�I*�O#S�Xhw% ���4�CSwc�Xx�i��x(\���Ҳ�j��ȹ^1���
�5,,����w@�9���1�8�%!!KΥ��j�Fr
-q�%�����!�:�_�F�W��)Sdɢo�9�������e�e�s	|��W��k����,�� ��̀	d�$t}��5��]Gk�����D�x���|Ȉ#w+�'�!++�OmP��ò�%����16�\�Wu����R���S9����0��Z;(����y|ͪfa�Yp#���\˹~�$ƗqdM:zzy�ڄ��WS����7cjkϓ��Xr��� 3u����G}�Ʈ�Q��x��ִ�tͅ��=����l���~�@�Lk1U|����GC� <��.-=�e˂���?e``��(ר���]�lvB6ݼߕ�M����rճD�q��jvߑ��!�7��(��T������ݳ8+I����	qꍖ={�����ft���*�qqq�x1$���8��r��EY��+��`{��:�:�q��&^Im������7���-.,���@+z��������t�+[�J�$��a���'wRT�BU�x�:.·w�&�S>�Ҥ�˷��kt�Y��N1㗅�/*�����K���9�g�����\c��Q�eEL�����M�g/0L�#I @�B��!j�OIr�Ww�������M���N��^
�#����h������I7�/��|r��w�L�<A�*~~
�YB^�͐��/G]�6�^�b�l7��ހ��&k/��Vn���b�uh\m0��4D)eO����[��&o�hyww���Rn4e�UW��xU���x�w��ˑ�%!E�G�� 0�`h��Z��XA�A�".�N�Yʓ��k8�tB���餴�a�s/眡9 ^0~��w�_�6��3F7+S���zr?�)���⓾�l�<A\��ek��g��Ţ�����Fm�]��0V���+����ԥ�5������gl3����HW��;7��9�). ���/�E|�);�f��#WUU�_Us�^���H�E�i=�n޺�T�IyM�r�����[�eg3::�����I�㫸!��%ෟ�(���"\���P�,���bZcT'�Ny� 0�8����7����O����Ʌ�,5�(���!`��ٳȶ����&*	R���ױu66�=��q���%�]�aE��a ��7�Nn�~��l��^p�]滇�b\��R��Fݥa���m��\w'���$/�} /�H�1ta���ج�f��O^l�5�|�^l�YS�\ t����@�cR;�Aoˠ��T�:ʚ�1O����--O,�����q�C����ݔ�S����SP����"q����a����~�F����TUV�ƒ��o� [��i�[@Bnpὥ�]��2�����X&Ld)S����,��/�5jи�+���Sa��--���\��qǉh!?���C�D��C�Qv�r��7��{M�[����7����.��s�n�̱jԨh��?���Aު�7t��3&���w�#� P蔶G"��@� �a�v\����_�(��"ۦ��>7g��аPW`�U-�`�]ܖ�R��"OKؽ�yX�.���L�w��z�|���o)F������5��-5�EFզ?qq�f���<1������ |b&����GiC���W q���
q������Y:�~?nk���hB�235���4�EȺ����0.��o���`@�}��$��quu��y� u�d�P0lѩ���'�1;�*r{�ې��w{z»x6��J8�����B����(TmC�	+$���I�ס����� 5�a^o@4z������5333����yy�p�3�zAƅ����d͏?��&���O��3�Z�G�[�Y��k\�-��Zs�Z�N���,)'k�b�Rz�毄�dPu��ٓ�
�8�"bA��$��	�>�%��i'CC��C��ۉ��� �DA�^�elll�+4΢}���' xV]A��j$���b��)u��-4#
�%���^s���U���*�5�E�j�7��fh;#�Τ۵ ю�)��m�=K^���-�h،����(�j�}����-�B���k�T�\�y���^�~�ݘ�m�O��!���2V��G�#�����W�I�M�B�d�+��E�p�M�.���^W�3~��n��D��dj���?:
M�Țȼ��Pʰ4j���_^.C�ۈpxP5�(� ��f�f;��.�d��SVV-=�	>� �H�@��W�7��D��:�4;9�6�󤘘�<"֢�Z�#�"{�����	���f�\�HY!I����������y� �,dl��
�@7i/-�,W���?&��pp�Ɓ([ �-;�w���d烇X�`�e}����P.�6�$�����.BJ�CI��@࿦"�-$GV���5*K���͚l��ic��_8;5��D�~��D!�=kћr���O�Nۑ"\�����7�����GmB�w�G���P�^��*�(��,۷C��GE[$	,��i���Ve� 	0j;�r������5���``N�0� ႁ�<�Z����D�N�iB�p�%�R�^;;�Hy�[��'7�SfV�҇�yڨ�*!UNQ�y�Ĭ�3hܳ�ewvv�@�nyz�y��/�y, Yʏ�t��n��
�����@\^C�Ӌu?pB���ID!;����܍������b�h�3;�l},�����F��Ƃ�'����(����BhZD��A���D��ᖁ����^��A�w7��mも8GCk�Z�g�q�^PXD����Ӣ��,v�����G�!Qÿ�t+�zv �sݸ^BRtS��.B�H\��+�L8s��a%W)��I!O�0����$ ����=Z�E�u>���9ȢI�aq_lEhl,�e���l02)�}.쯿�"�\yBE���3�H��ʲ>n�0�a^(�ښ�h�̶�R<�1�v*�.�#E`�
�9'׋1Q�p� Ty+����Y���Ť?�Mc|��ڊs�Д�ɔ�ag!�S Ehs��� �	�����ؼ9"*�S������CD����m&�g��Ͱnjg�^����6���yӄ���ڹ�&]%}��O�HJP��W�������:��[��]�*��p�^��a��B��U��'=�k�^^KVڹz�L��>N�s�R�:$3-qf�a����ؚ����
l8��t��$�~�4n&x�̸����������;�HJn�d�����_�˫��O���653�DK��B�	y��͛n�PfoμW�1�d]�L�{������U�zzhi�b���|cpA��7�O-1 ���/υ�7~eQ�KJ�L��A.x/p*ـ��o�k:fAL�'�����d>az���_��
p�4&�L����׍�࠱��.��S]�A��J^6��P�]��4����~���YBY���˗!{B������A0�|k�<��Md��틻�!�i��	a2�[�����K��K��j�s�!�F�3yS�@�[:��y��9{ԯ��Bl��7멐�l3�B��_�>ыI��W[�j҅�F������,6���4i֕�oa�e�s��Z�����օ����ߵ^|RS��E��8�o=�ɵ�&�lVW_�%�SJ�����%�CVRJ�3�.a�j ����)�������	�� eO	����.[L�S,B�Z�9��>݃,�5����ӳ�F�lS�9�/����ޛ
�k`p����t��i�	~|�ۓ���(�J
/[Ԛ����P �<� �ŁB�DO9�U��׃«�Yy�{v�G�r?�K�ý!>��� [t�|���( �-"##�{�F�a�h/*a��Gi77�pj�o�/����Cv���>����������;����S�����k��D�����`��e�4x�y!��3�����Pг�v�_��D|$rr����4�ir�HS������;uOI$��'��č{N��g��v-ҷ�
���fgvJ�l��f;�t�G{�ns[y�:l��+�&�~Z���~�:�����ނ:��إ��D��"�wڜ\AcM�VT���o�� {tK�?ioH5$�p�����{K#�&�X�������fo 6�Á!�9�����t7���W=��+"�^�����p�1�����	e�[`�~!�5�߸'�vm�a��;Ӈ��Nn��#e͐�\ٺt�֨����_B�ۏ�>ccc���{���W���b�#AP9|����4�?����٥Pg��)�d s�g�"���v�>��M�o|�����/>>�v�"�8B|�Kym��*K
�j�)~�;L$�<:0e�󬰰���x{U1.,`^)&�����1�>Pboo�-y$������Ե� ��<���(���s~� tZ]�ABF�C_����O}d��,{!�\6�����!�]�^f5j�,:�������H0��"�wKE�,��wo=G0�����F�[��+/>F~9?B�PPP`�i��0�֭�?at6&&��޽{��D�� ���؃��F����|��w�D�����S�4���4s;��g�����_dU�:�1Vp����D�3r�/E>U6�<6ߪ>�!��a'�+�U���T�&� ����Y@@Ey9��0�|����� ?Sè�)�b�}2�6�"�o�q�b�~� ^Qm\q^0\������n�=��p����T�5MM����A����<<&�l�^[[�Lh	�o{wP9�`WIH	�`n��f��x?ga�`l7��c�!��+(��R�A<���Fq�Q�`pk���OL�n��r�x���uȫxf�جg�O֪�qH���l"IP!�ߐ��,�~�T'vAgvrH)^Kz��ا��HY\��Kb~
R�����O5��^B`����=�|)b��è�T������&�4?
���%,H����/E�����)y2+����x����D,u�3@^M�L^�0�=R�
�;
L���'���oH��Q�o�q�@�sI0�����n��r��&�	��@�0Q���4Y������xw��9�/R>b���3��_<�=��HoTl'�N[x9u�<#p������>Aj�N��_�S@��W���v���<�����D�^��
�1�_b�?���$텪�Rg��b�� ����!��=>�UңL�LO�Q���_6XEk3�J�V�����&&&�����oU��cV-N��cU�?�a0\�Gyno&�!o���czv˝�A4Z`s�Y��旇�ώE}ݯ�F'N?��K,�%I����Z�C?�qx��R6npݕO�F�W����?jѼ�
��8��e` ʄ�;�~$�dAU`���l��>�,P%м������׽W�S#�$���H[����羢@���|N`���`CJ��y������U��V��U�t[��y�c�pT�Ƥ��D,��غ�С$��Eqd �Ԗ�D\��޺�)��v�lllf��D��6��a�����VC�嫄K���v��X���3�Px�Y,H� �U��⩥3�@�i��"Yd i@D1���G��w =s��
ѣ{�]�jR?�J@r�]�Kl�U}��m(b�s|��XlG_p���駿Y��5�l��]�3���oZ��'�4:�@y�Pk�<��i=֓��xwŧq�����%�JĎ�Y��X��G���3�r��J��.��/ y��B2>Q���v���p
���:��S�_lH�οU�&��N��fVo`���n�ϫW�p},$|�tSiIUMM�Z�ɿ�����.]4
�.�;���+P�!L�A���B�C>"���R��h��q�P'�}[�	MR����Y�� ���>x)�Č��At��Kn!�q������5�G@����p|ρ\C�1����,���;�531�0C����p�0��fL)�8'%%e>Ф
=Z��#�^� �	�g-��T.�{�����d-�D�"�2 �lOY��"�0v�������d��h�]�iRn�9��k��\�&L�y�?���f
�\����ʪ���Uʹm�v����vN�<yY1oJ�v����-T�h�VJ��%h��ޞ�޴A�c"2��%7�+���ӊ����ۯ�=	�6)d��c��&��"�B�����#�T��ROT40�222����/{;˒��gjKn4�A���|�͠�M�Z�jk�qE�G���� 0��=y��jbLMM��^/���1�|6����!~RA��xG��Dnh
��(�@x�TZVSS2���[}rW����aFډ� �%�l^{�6EPI�F�'�H~؉�PJL���o�h���|�8	����sD�,� i�6gcc�)���P$�P��I�yMڹj�̧����|�f^J?9�sE9A���`�@O����o�>��yyx�b��b�7���m۶�o���f&��&p�U����O�O�4�)�@�����d3!�@@����4�t!��jT}���p6�
�Q���$
��OdC�F�`�e� �>?9"��)���
�7�yTP+ ��V����n} �G��Bŭ�1=Y֙`]����.,l�Y#h��s�QMooo�Tcmԥ�Lđ�6�al�Yq)�� �`^�P�?FR����^?�PZQ�Ѷ���}�.�rU�!S�o�,��|
dW}�em�����q��H����ʤ��V���
��y�" c�p������3\[b<d�2�A�ݾ�8M)����>���K25���-�+��,�;��؅����T�8cc�;?����~q8��\�x���Sȴ[�LZr=JB��.tv��ܔ�}���E|�S��H����f�ׅTVW����Z��[�6i!���ë��p�B��.���鯯/���j=z�����R6�w��Hun���\�=��X�
V�폌�.p�6�b��R���c��7LSi��	�dJ�Y�|�/>]��p���SD$ip�W��I=ڑ7Ԗ�vao9��q��dd8�1<<<�QRb��c�Dtt43y�Sٜ�;/d��9�@E"6f <���s��m�st��O�w�����	2��V.���� K�mO�7�56k��<����W��!Q\�E������L�w��	�����#�.�h�b��8�!>�'ۉ�Ɨ��n�����3 Ԏ� �@� g1s��\�>�>?�=/�n��-�z��'s�w��&]����R�I� Q{w:��@@b�X����i�jbe�tK𚇡֜�o��><��K�C�-89q>�x�c)v�������<�O��o(�H2�*B�:��hW�JG"z
�rqad˯���
��8��g����$�FGl8�h��R�$�F����y��ā<r�!�0 ?x�j�z a�o����@��c��F�<��OVS�#�%Z#�EPK�\L�t/V�����#���ő}�3�qf����C"O �	����5 �WJ�u�J���D@I���t�D��a��y�S�Ne{Ǿ��!нʴ���)�K�I��G9zo��W�-<�]�/yK7��{֋�)	>~vWȤ����Uk/q{77u�JjL�r w�L�06<i�@�Q.��K�Uf�_�t���+'��Sa8�e�\⃮z�]D��g5^�3�y�l��8�S]DǑN�6�t�@����^�k0c�3�i��#^������O��N4�X�R�f7��@��Px���VEA\#"�{lԧ -hP�UsM��l��mhr,p}���,��=�>�N���'9��(��$dV�ӫn�aV?��_װ��v�7�.4/$�����	�~R3~mV��UĎ��ԨUG���d�2ż��>,=]D���en���92�4�GP�����mO�۷?�E?ĂlSN�/zvLo�O}^S�zH-��8G�����Y4����q��.+6�0�_�h���
@���c���H�A�Y��!6���"��HM��&�~"�s
�� -j3�LԬ{�q˻����Ǯ�@�0\�Ϡ�����!ߛ'h�QAA���*�d� �F�#8+�y)���NN�o���� �I7h���Xz��V�Aќ���fͅ'}\�zյX��& �Z^�/vٺ
R�e��\����`�NT��zl;|�o�	��t����K'�7�S7
��ޜq��0�/���i2@لX�*� `c~S�M0(�K���x9`i��
`,��X�\]�>��Ԯ�����m@"}��F�JJ@
8�gq�1h%��?�(�ع"��i'�ֳ]�!�?�W;��%h���^t`� ��1�],�����qJ	r�����H�>_� ��<t���_��͋( '���y��=W�����!�m)�y!�y!Z@K���9���g�l�
�C�I�5j#F�9��q!pK����f�t�sF,PK<����]f��yr2s�Jf�U~����m�S�L��o�+j�=���d��ma�	��ܞB��B����z��^�%]PP��usyMӎ�%����vf��APǖ��s�|߂�C��x��=��t@O��:�kY��)L�0�x	���o�fpQ�����}.k�U���D(pg�THB�'4�T��-����� �q��6�w����)-V^�W"��|�1������x/C��	r4`�����^�\�wI̺���von�<���6"�	��ː^@f�N��`p�bQQ�UbM�f�#<W��,oNw����s�AF(~��p	��ϑ����;u�N��^�u% U#�|:]�A��m��!0'=~�U\\�5g�^�10��� O�k����P�^���1ș~�H���X4���Z��5۹n�*Uh��Y�e�c^�QJ���{��RǪ�M��F���WG+WTW_1e��I�������q+R5%�I�s�Y%V#ͅ��K���Grc���ZGr(@'2/�Б:�X\�[�����M���8�%DN� ������9��O�AD�W�*�j��vs�XWI���=ni2�,���������|��a�@䍍�����L\���<��J8�= �:r��@��?������3����1����z�������,[^GF�M��.��5�G��������v�k1�C/]���ZgkApiiF�����W�g$�<�K��8�E��X��\�t�~�Q��):0�8��'��H�~��#�]vX�S6�����\����/���逵��b�&^�sL���2��!4�cѢ'�h;0�^]����x�I2�cйZ�o��O�S�Ĭv��!V���m	�}0�g�����^�*�@f�A)"�~����X�6]]]��w��M:ρ6Y3)bi~��.�[�wcmt����E4@���qڝ[x��:!�NaA���_�*���3j�g]���r�*�a{���I%1s� �\~GL��c2�)� @��-5ʻH`P�qd�� 낂���E�L��}��W		𿙳�c9�UA/B����3຀`������A�+Wn��DFF�^VUm�?��	��U%%�����i���^ 
1Ԧ[܍�ٞ��@� �Ԭ������g���:ǂw�Y1����6y� ��5����]#x�~��A	��K-���P��t]}��t_�Ns��ρ�|�JV�0�D�����@�O������6��M�J�DP7��'�B�k�Q����Q��H �_�Q1�@GVU�;�ׁD���:	'�\�G�(�^�O9�~��D<	j^�|đ[�����j#0���U����ٌ�P�!0������eho�eHp���y�j����~C�Z�q�� @s /�7�.s�'k�kHOK����~{5��X�g?	�`�4~�� ,�']�l��q!(m��~꺪��g���<�����ׯϜ?_t7Z���
z7�Cڸ���d4멯/s���d��4k��	�֣˷;8������<�Ĳ��g>vg�;�:��a���2�.�=����#�˗3;��E�/\�|���
'� ��w&�QVq۔�j����Z����S�tQ�N���׎��y�3h�@\���d���v4�˃�n�]�߆�?s��Z��g�(��*��?��ϐ���7�oKA� ��Ѿ���#8�0~|Sf7[���,�~o���w,m�QCY��(E��g�����FG`J[c��4v�1m�5+U)tN(��|��֋�ڛ��P�����ձ���*'��h�<�Y�G��/�ߔ)�(�G��Wb�{����3�j�Ӵ�YRt$�aЗ���T5�h�$[�^�}���7�f�TY�eo#8�h��%.�K�t�9ٴR�1��x����z���9�a/��GM��3�9�؊���+�8�V/?#)Q�9"�S���D"��X~�t}���q<�C%*������(�f:������MOOo����6��/�T��JKKn";�m�Z�����3�t���~�J4n\�X>�	�!7���p�r��$.�L��u�k ]�VwP=p�'
!�������H�:9>�w=U���G�l|�I;�oY�&�^;�����ˍ���� ^��i�v���7��`0�l�XT��!@XD�f�8�m�0�Mu�x�ML�@uZ���Z��C8�Șiܯ���3jB��TM���b�V��I;�,�ö����L��c��uc3Z��%@�C�TL�
�P�Ĥ��<ΐU6��ĹҰ�H��{͗�!���\��љ���S8��r怣�Y�P=$
��7{V;�9B������ t����C��s=��~��&z*�l�p	�#��'Xv����^���'6cS�9@�Lk3���9V����<$&�n7Z&>�}��.B�0��W":r.�1���F��"՘;�FˤLȳS���h'�NՖ����>ק~��:#7��8�Y�|�#��؏'��S�C��n�3u�AYV�C�&��v/�N L���뛙ͺ��PjÅ���W�&�@"�O~��j<�~��s�)#����!/<7�6�@}��-����� �M� ��Y]W�,d���nc�:C��@s #s5�����M�M0�	ҳg�Q�PW����ꍌXs�[�v��L����e�3�������"�`����ٿ�ĥ���|�^KSU�7N�Z���5((�)����?�0��moWF��'?b������%��$n�q+�z����C<P���e�õ�����}��F�~)��
$<5�ŋ�O�91�+�jA ��~�Ձ��"�l���\���:d���Zl`/�����/������޳����@�+����\��`1�_�̄�pc}5�AC��爙�m���6���i��/cx��is�j}��ky���)	!�a-x�$ԋ��k>�z��%j��ުS:4�pB%k�� "!!aiuei:~�&LEeOG�ZX0��� ���_��@�<yb���G����!��&b��awf���X���܊S��S�b��KR��)� T�x"���dTF� �>b{�M����֡ͽ$R�E�H�k�q];<
$�	��e�/i��X�=�kq�^Zs�����_�3�-f3���m^뺝l ;@�/���~���w��xrvD�sy�ZG�;�&&& ![�{]ʇ�К1�	+�~�fD̘���藪�$����\�)��?��Q��5(j�K�!�n�i�p-���ˁ��ƥ�S#]n�S�<~��͎�v��
��¸����s�b����9}r����_#o��YV��/�=� @��b�K1��4Ϩ����aI2�.�ʄL���~�.p��9nj`~.���_`Y�`���^�a.v��YX޺0td�)�1\7N�	�~�5����0eO+Ld7{i�z�+�;�4.��"�e\T�ub�o��������)�=�ů��E���`�����9����p�}��@�sy�'�=���;]$f���f�(��|��)��T�
�_��m�#�v<�ي���aX���O�P&T�,?M�g��.8�n`�?{D���cf?��.��y��Pw���_�S�-���U�C�<��M3��؁��o&�S��l�\�������|��� 
P&�R�@���`xv��9�L�^�j��4��kl���X��'��tEFs��]W�dv#�ƒ�E����C�q
�>$��������y��.�[���s/�zJ����w?|	i�ܶ�G=T�/�~/hQG@��ʂG�ϞH�l����?
� uCX�C@>�����H8����mm�w~X���Q�	��o���f,G�փ�����8ÁgS��뮀�Re��!wʤ*U���U�d�'�~����q���(�<���7����g�j�[�N����NX��
�}�����t���z�M�6nz�f�|��2�x<�!�EKϨ���]\�ݵ����j�5\d`/@���Æ���A7Qkk3fPq6�f�C}�ϡ��B�/C�G��:����H�����yj>�\�������
�f��C�,qf���P=N�^)?��@1SPy,k����i��CJ)��:]�	�}��%I�aLS�nZyU2�^c��k�/���}��������J�P���t�_�{���\mv�]���K�rgY����(��R��H{X|g��2�N�K@jXW���XI�	n,�n��������zf_>u^�}bN3�G����J�����20���O��l!����ƃt7ˊntww���xƐ3���{..2���V������^��W~i��1*�����?~\.c�ӌ����}<�8H�Edd����w:�1�}��ܾ��#�bﱟ��EB� n��%�bTC|��Ѣ�}nf"��]��+��8'������fև�K���U�pch$d^�UD�>q%i"���P�����}��pHto��C��\�/�鯫n�w�Z11��JTN�|�uc�#u��/.E>��ˢ�����a�!p4��#�4p8�e��l3�Ɍ',LOO{�S��ٗ�\�y�\f���]��x�Uz��+t�z����)1j��Цd2�\���i��v cπ�w�Y��"�J����
7�М.hλ����|���DϖP�����������#��� 0`�'+I�?����1?���nsQ�l�[�W3��y� ��߸q�l��#}�$(ˎqMʶm���R�������Y�mR�vp�ioN���}9����ǫW�~����p�8��ˡ�=\#�3����Ƈ����Kԓ����2ǉ��:ũ�N��}�xN�ߜ�V�l�q6��5��Ά�U���]$>8�����s��mLa6e������ 
�����)�۳g����c�aX�9٬pvv�3�)�mk㵩����{�Q&-���LK�g�ka�3 δ��R#��BT��T�o�b���4���@��-�_�1E�g����w-��;��9jZ�N�F��e>l�b�?�Vw���f}�9 ��=�Q��3ý���Y��+&^��F'7���|K��\	���Z>ˠ�*άn{�����CY�ǻk�|�o��2���R�_B����E`t���w������]�O� ���]�d��+�W�pZ�3�I���#d�������W�0� �^��ō
�z£3���b�������K��0�[��w���}�����W��:��7���8�5#�3�n���GO8e�X�ۍiǶ�P���#'N�H�ԖPn� =����0$����o���Ϝ��>�#���\%�"�<���T��׊	%�7�������T�UWo-**
_��� �1333�a����Qn2��GC����X)�;w�|��EԶ�<�^����ge�����b��<����<��ێ�'QWF�5뭌�̓�߄GEFU���V7t���1����a�UR�Qז��͎'���b?,$�d�8�hǈ' =~���[��5�J1�)?R��,@�+�"�UMS�ה:�Gj�O�x��|�n��x�i"�O��b����n2?�=,*�b�f�}�]0�3���f�r*�Ң�30��LO.�����������:�t��OF�=����8���s[�v�/8?_] ��ҙ�hl�<#Z]YɄŵ�
iii�x��� ����?�)f}Wz�D�^a�*2uNtn�b蛦�w�20E�DU�N����-x�Nî�����N�lV�b����啨S��qP$�r�gZ�������� ��/��il��n2:1��׊�>��[{"BA8���l<l�aVVV����[���Ш�����y����	�A�@1��Q�M�RF� ��J�6<_�zv5����	��E���~� ��@��P[�,(8	�U��	���Err��N��i��R0w������ˊmQ���|�ÿ��u���se��©ٍUY��MȔ\�j�,2q��z������O�C=��m'g;��K����]Ij��S<9]��Σs�*:�h��/��H]��N��v�P���ÍKH����R'����9�Jo�8a֫Py+����J�(^R?��g��Km���=D]��i�wK�����=��BMx�iݺuq��'�}�w,$��2>*{|�o�n*+��y!𾿿?��^3�>�t�F��N����t�q���K��oH��ܸ\�0@�Qg�?��E�盪[=҅{VX\�'��)[�I�[c����r����]�^?4T�l���-����>��L�Х��c��:��J�ˤ[Uo�z���w&�rܘ۾�i��ֲB��"JlL�������t��GT�z�.`!���x��I�m�9�wRn�ō��QWN�����L�޽y��A*����q�n��VT��C�\h��f�!b��'��!r�"mGݨ��7;��3�:ϯF��
��d�a,�$PĂ�{�F�7�O�RMt���渭�[F��y��VP~xf�	 ��{St�u.�ݼy���z��v<)p��QZnE�7� ����A;�����eJ�=z0%���8�����������cc=���9�Y~��]��@�����{w��IWq�ؖ���y����H>�	��	���ު(̊W����Xu�u��?oK�@�Jʚ�9 �w0���W��ek(�}㼼�Zx�3�s�n���_ܷ��w����ϟ�X�K�������U�`a�S{H&�''|�_I<|H=K��իxH�E	���Snge�%��g�]���R�;���K�Q˴N=z&*l��w����׵��B����f;5�O�x^0��]ӫ����oRX~lY
���p��Q��'Oᰜ�@~c���G�wv ��9k�D��@�>	�K#<4�A�C@���-<��q(R֎�#NM����2J�����fx�4�-�Hr�����S.��T3Ѯ�y���K�>�zeB�&�g"��0�	lO�=z��)MM̓J��$������^�O��o����2aݺ�1��?[��Uu����C�%P���p�����G�3�B1e�?0�a^^� 0����o=�J�Zu��ƻ��H=Dp[խ1�6���\\����}i��J�g~܃?�p���s�#�2g=Z���� ,�q��@����BɒkVPٽ�!�J%z�K����ȴ�
{/wR飝���?����w����]��*W����U���w����]��V�8_�V�����A����׎$�OLW����ΩǤ��4�+�61P��������$�_j��K_��@�ܕ��-ZMG������w��+�]���
y���!\����+�]��
W�������w��?Vh���@zL_����=a��pqպ�߈"��M�-��IwB~�����G�p�o]߉�)}���1i��� PK   (_�X��D>  ?>  /   images/61ab5d34-94e9-4496-9157-f8e280b3269a.png?>���PNG

   IHDR   d   �   (�-F   	pHYs  ��  �����   tEXtSoftware www.inkscape.org��<  =�IDATx��}x�u�?3��ŢW�;ER%QT�:-Q�r��{�{lŶ�����;Q���ʲ;J,ٲ��%J�D�)���lߙy�3�X� � Rrx���3;3���Ϲ�����6Y�H���K��W�৯� �� M�m[�/���%���q�?�o\W�eeAܳw �n��-�Ć�����߄������x�=�]�q�N�<,|�
�ǎ^ܱ��H���P���ڃ�T��>�����R���`wW#㺤.���_�i�}^U���룿oD����?Z�C}1lk���4>�6���˱q� ��B'.^P�Ｅ^��?f�}�(j�eM9n{�	[[G��˪q��R�b{݁SʲqaM>��H��6 a����m�l.JJ'W/*�W���gj�ֶ(���Q�0zQ��T:GS��LbOw����͈���{����rܷߺ�߹��!�:2��܃=�yZ���,Ë�a������\���X+�m
��7�"����>�'���a���c�o�`4��ҧ&��2�no.�y]5�ws=��a���](Т��>��>75���o���\��է���������a��"L��B �[F��&�z��De�$�f`���\|��E��CMH�l��YA�r}:��Z|���jB�俄+CB�y!tE�1�?߱BQ�uK
q��-YC�5�i�]�.�h�U�|����P+H�_����&�;�� ?A���J�z�
|��fv��t6�ޟ�ׄ�$?�����������|��||c�Ɵ�=�5����|h4qW�*���6�qmF	���G���/ .綍��W��	!��en��6�]y;p]�>���<]����S��ѵ�������DU� ����s02�C��g-|���p˹e�������g!l~a�p����$��;+;q�M�CqYZ������Q��ޥ�]}
��l�[VUa�5�nx��!�m�{��p������0ޟ�7\}��}£�����ۼ�/����й�7�&\}ӧQ>o!ښw!��_H���~]8���y	oY^����,�� v�|?��6�߬w�+O���T�bx�9�t�z�u���EFP��O0��
�_������`+�]����	̫Y�ζ(|�5�Gె�����꺕���� ���W���/nT���#��G|f۲B��@"y�u�W_�Ҋ:un��uX��,�ۊ&}|B��ZKs��z��#�d[��f�ڷ�!te"�5�i�XTQ�kެ�)(����Ê֍��_M�[��ҳ.BE�bu��Ek�x�
,}��Z��F1,�uK?��P���7aϞ���GԨ i��{��4+/� �c ����ވ�ͿV N	2`�X�&,Yv��P�"З,=˷6a��P��h k.܀��buݚ��������t��f1��Den4<4�|<��e�sK�MJ8"ajB}�n��&Yjʄ}�lg�	yV<C2W��	ʳ|���,[�/�t�5���J]�-}
p�Ȩ�?v��K�L��H��5!�%!b*� �[0֧���aZT�p��g�}�w�)���F2���&�	d�4&���G۴ �Z�q��'��W����hܻ;ۇ��Z(Tm�T,��Q/'�b�3w��7��Ϗ][6b[�Vc!*B:bb}JV�~���pɵ�����a�y���a�XoGGLl�Va��G�W�QQj�����҅��:4y>��H��X��=�̔pf>vo} ���q�,KK�t�#�Jl
���;�K�Gx�OD����y����i�}�ī�Y��� 
6�Vqdk�v�j<��[�%8��/z%�����)�K^��8�AA��2�%��,y`$ea$n���[/%�+q��Pd<�6�%7`��ÿ�X���d�ȽG���|$;Dw�w7(E����(��"�����&���k�Ϣעg�,<p"����ǖ��V�����}Q���`�Ǹ�^A��:�B<��]f�ym5޲���	���[î~�fbj>�_�,'�N��н��El=����w"f��OEW���y�R����M�g�Z4���[^B����Rע9Y��^=�?�_x����FF���o'W�$/��ɸ~��C��,��|�)|�YQ�w�c���w_�I�u¼)D� �b��-�1,H��#-b�/��n�}m�I�\e��
����S1-��b���w�+���؛�J~GL�[]�O]T����_��_�\�7E,�K�"GP����u���	�*���u���O����5x�X��P�Y'\��w,�Ϸ�� G�/�Y���_F�F��Tb*,}�uy�xy5n���]<���*|��P�f1Ɠ"�Đ���ը-��C�k��lӻq��A�JhWq�޾���bp������B1�I��s?|�B\/�m8�(+[�U���v1��"f1mn��o�P�va�4��u�ů 2����J) ��-E�x|uѢ����}Gā��֍G��7/ă�D���|4������GZ���m��lX��pRܱ�/�'���R������o߿D8t�O��hRN�m=��1d�C��>�����m6cT�r�b��Ou�5�h�i
��kg/~(�mȟ=2�F��P�`,%�u�~w���qyM9M���A��K���k�*/�Q�~�S�hPy��x]����hJ]IXʳ'G�	�}
!�A���^�����I��}���#quۏ�u���!E�v�u��I�>�%p3�����q�Kyݾ�(>p�a�����$�bB ��t�1-���e�Fz��!�y���`�PSf��߼�|C-���^�����Lѧ6�gO$��p��g��rC� ��>Ǯ#a��)���<���I8�"=��S�C++��.۟��Ag1�l�<|��u�'a1C�Oڦ��3mn����Z!TJI�	�Ol41����&k�i�7�"�27�sK�	�ØM��o&����/�;��9n
!I[Ǌ�!|��&�-��@���0O2C��M����芕�P��h6�q��;ѧ>����o
ꎃG�9���>�rs���4)�N� 	�\��W'ě�g�6�R�ki���k��I<�>��ӌ��ަ�(N�l��(,Y
� ���JA�S��?��]�M	��u`�у�f9V}�nV�b�(�K�c���O-��<�Z����Tr1��7���u��4�P?�s�1fF�4��V�P]~nB99j�9�"�D\�4�g�jB���p�h�|�BL_/�z?L1<�i�>�!31� �TH}ک^��Q����S>h2';'�?��L���RB�<3�^|6M!��-�G�w��<�'0�8Y]�|�DW�1Rם�&V����|�Zl�1�r�E�"�r��O�Y?��/�)��O>s�
rst�KnAϊ����969c^��]��(ׇ��a��\}�C��
!\n����H�}�twU.�&�\�^C;�<"@��F��"����tw�'sޱ�#N��g.9�f��@�f�����!������̜T݇���c"K��D�1n��y�5�$��i�N�Q;��=�S��^I�R(��Wˮ�4��J��u�=Iy�֗��M87E���644�Dr)#'cٵq�:��4�"���7d���K�:��2�! 9I�h�̈́�x�_���>+��r�ײD,������Y&S>W�O�Vݸ¿���*������9�"�%�){*���x�g@��Y��/��c��wc�]���H&x�;ߊ��K���� �^W��'k{q�]w�A��/++ŵ��>�9���5c'��p�9/R@%�n�0������s�0����AH�7.���?�H$� LĿ�������@_��=����J�Al��B���X]Bii	��[P�O O�*WK�di!P9��Dm���E\͛��d?a; ��,6�#�IB!8i�K��;��'Ї�s�g6<����E��]
��s�X*��v�8���\|��O�8h`0Ǔ[��x�I�\�
����^���$�`$U��@}�J���̿��yf��L��4���k����-7Ll|������h�r]<1RRf*�%C�`�I,��c��DLh��-�����iCi�����[<�қ1�v}����n��⊍ruOo_�o��$#z�D��'%��]V� b��!>)*�� Em� ���Y���1T�ּ1}�eSLL��1�}��]�cV�fFyY��5*V�Z��#��(��8,��!�J;P��t�ir�7�?	��.��".bӢ�5>)(�[�<7�坐C<��	A/X>��"�|�䖧2f�Ī�Y������2���C���˗�I5�e�I�,���>��#ibT�S6f�\�S��0��(�8��z��N��23m����K�8S�*�R�H�$(��d�>$������"�D��V�Àf�H����s�z�ODD�^�-P�)'l�G���R`pUy)"9�hL�)�ז5�ׇq�����P0�E�cǠ������&�p�,�nj*�8{b���ߜ�^�#� ���ڢj�n���◝�t	�Gr0��f)c~�@���}~3^���8f�����T\�zi�>�{�,+Kt�I�Q�������\�b�����񛿄����x0�=X�>�*�G�>�E!���Q��ڑ4�D))$�� ��ea|��w"�`������Ư��ʰo�L|O�?�����9C��@;�'����.�}Ǆ���b~]bb�����N&�J��ʠ[��!~���A�rJV��1���B�WU�$FOw�*�p�D��.'�ru�v~���G�1|��a�~d+�Ǭ,z�@��á*�~�|I����q�?�6���gPG�U�����)*).�֣�%3$�L�_���2�T�oSot!��B3�O�������Z�"ĺ�
9��
�D��c�L?%C���P��ʪą@��Y�ɢ�BS�_��d��sޜ���A�pL��1G��r����Ю��;�E(h�az�3�l�)�����$g ��j�V:Ru�<!2�/{c6�z��%���?��0D�O�~����$���4r�B�AX�Ō���+͘p��N�����a�ј9M�n1%�Z��a�f����b�-�5`�Y�v� ;�5a�l�oj {�?�H���9^������sވx���8v|P����Б�*��/~�Z��!;2]�P�$�I�� J������?��ؙ�"�!�8��ԩ�h��˜����b�מ2�=��Ԧ����̞d���B9/��D8��?֯_�b�!ñ6��5����� FlACc���L�k�C{�Y��p4h^��̇���'�N�,����.cbIk�U*�G�`^n���m&�A���ƺ^9�'�<[S�V��D6��>P3�{�W-���@ ��������B��v���9�^z�c�D
�ΰ�qg�o�ch�� ����	(?dCQ=���xC�B̻��S��yQ��2-��jq}�����"8��RN,'9��{tM���oR'�Q�P��a4Z%X.��^����kUb�ރb�3ڕa����#�eH�8'��9�B6Mž:�W��+zȱ:�C�DpU�[�@�����VN��m|m�h:�'�Чh���d�=��c�4��v��$�M9�h�Zu���\�Ԉ��/��M�b��S�Q��pj�5�R�Q/T�/��ADcLr� �T�6L��'SɄ_y���3��t�$�]i�PGܳoV��u7�W�s�38��rǮ�������}�oN��C�·6w��Zx���l���zm�pF���D���>q�"f=��\<l.��<�I��s�|�p��X�<��ʩ���4���F$D�)+����,�O����1�Hg� �χ=�Pk��Β	z-���M��訍_�T���:�e?�]I���x#@�S����6��g�JS���N��G���H�8Q�=a�n�������"�����m:���t˩5�(i�`��b�%!�X���Z`~�K=�ŵ���k��R�5�b�7����F {~É>}�gڔg�=#�K��&�I�H����BW���ocK��2a2%�8�0TpAA߸��ԕ+��VC� ��y����tI��n��m�c��z��n��*�H庖�Ѣ�]A�_�|��+?����=��+)�,#��ǅ�ˌ8�����cݝ_6�)l�Ϳ9����n������:���@�>)�s�8��`4�k� ����'B
w���R_�aw����2|z^����ӥ�i�p_�kꃂ�E��K�j�Εa��� ,��U����w��]��PQQ�?�)|�8�������Q����-�s����yJ���m�����&��\K$�tA�%�㐑n� >r�"�d�&50�YV]GU-�.�NUO,�,�5P�V,LS�X�GI.�B#$JC>Ya��ExA=����˔:�A?�+K����8��b5�ŕ���>~�1�.fm�p4�$��&��b�gOmc$iT��MmL=�/:�}�#2��	�'BGR��WL~�`�D�<V�|;<$@�ca�9GC1��;��:���z��dO"+>����=τ��^�F�Z����>��;�o�o�0�O��������v�����&��w�����D�ﮰ�SÝ�\����Z_$�O�߄��Ѵ����΃�zƠ�ht8z�-��;�9�vv������X\��/��	��϶��av|���l�q���;�Z��pT�S3H��Q��4Co�v�s�4��}����Ǖ��/����a�M�'�$�)=�$~(X%��hW{�a�)od ���\����ҏp��c�n:!^��Z��s*u�hg�0���-�&b���qaNu��9�\��
�{���Ԇ�i3k�ge���j<�,z
�?�RW��y�*Kh��j��A�����8�-�o*y�,�����\R��s�)d���ˢ
��֧~|C�
��3��XW$�����Y	���7���}��(
jxZ8�p�`��Ѥ�m��V���Z������+D���b��AΞK}���ۈ$m������f�����5����)�����j/
īX-�a4aco���i�Q�4��*�q��H��"b�K>��L��yȑAK))C�b��2�~�s������d ~�=tRq�{4��S�M41�n2O%��{�L��&�s�EE:�_�����E��g	#���L�	�.$qϵaC�!pk��6����zC=|(ncG��t���R��s��X���y�e�AQrHwvD�v�X�q���ɅE�mn���s����AT��{��ykX;�=�gy���s��cخ
j4T�bs���H/�O�]�(��2]Z��&��Ԍ��-:���	Ǻ"R�%D�&�!�/�)�gT ��!����&��z�==��=`_�D�ʪr�YGGt��q8	81�����7�wb}e�e�Z�h�B��	|���?��%U��/Oq��rϕI���-)4�^-DMvOJ�ab��a|�r���C��j-Q���E�g�m*����/��a�r����]A}��HSz��A���(\A��ȡ�!�A���}x�1��;��P""O��C��8�T��.�=�!���,�(s8e�tB��O0�rv��L��?���m���u7�W�De�t����~+��� ���:�Ƣy�1�i��=���z��8U�v�ݏ�<��o[�J���P���w⎧~���G�kQt�`yr�����PW�T'��Y`D�3�2A�N�Q<]\#��d��VS��Ǵb���m�	�u��y��*!��4���U�w��8r�D������h��9 s�l/|G�O��ǯ	�>�K��2�x�m�{2�E�I��w��&XPU��V�1'j^���M�5u�C�t�vFhJ���7��v�O�V=�B��WҎ	PfWH=Uʋ�pѰ��
Ȫ�E��!�4�ISe:��@�ꛓi:���8��@ �J_�	�����g3�v��椒2�<��we�݉c���ZR��[e��jqi
�@wa��h
�)��$w�j���Y�s�C@o�J��J��r�;�˰4�:s�rm�ǚ���4l��N����UY^.�k�����\g��)�U_A~��,Q\���҈��	`ѢE�$�R���=�d���k�z��\�%�O`�h��Ԝm;<��mV7��� ��v�U���ը^yeV[Jq]qI).���*,�1��9&T���q�57�yN��mC0;R����I��g��R���q��KǛF`��QYQ]�7��3J����"Y�����#l�<Vxм���Nۮ�d��w$���BZ�/]D�?I_����z�櫉�N���'��}X��G[=17�I�kb���Q�%�4c�]�m���e���H����h���6�=����f�r�U�or�{�e�!1��Cfڴc�L�[��Ox�v��NQ��SiDؙǎQsf#�S��:c:x����{�������:ӎߴ����9Ӳo�:$�!�BNe��DV:�z�C�����0�������v<�׳�� �7o��t��K3� �4�t+C�x�"��Xy#5o�|6��,�{��O�R��Jr4�.�Fj�AM-����A
�ׁ�K*cJ�znL!������m���v��F-�<{�aym<�80�N���eN�=�[���"�By��z=��ziF\�~��ě�j�/3j&�YNM�xJ�O�RW���:��L����U�kX/�G�^WU���r�d"�y�Id����c�Z;���2�
?�}p��9HL�p�'���:��Wj�^��\7��d2 �5����
a�SEH�%BXL��k�f"��D��T�DdqAhe��2+�I�Mgc�y�R΂?�yU��i��^�3D�v8	m���b�H$	�CnZ�S����'�%* ڸ���!��T,*�r�T�~�F!��)Lv9�t��\Q<�LW��ϴ���^<j�A ESxhR�\0��e����1S��~����9A��V.���uRr��iX)�&u1�Z#��)�p�ٹƴ�NE�24�u��
'͓ ��+��3�:l���C�O��y�7ݖ�D=qs&�8AV]Ѳ"Փh��/�F��I�-(d*��-m&��8��:��I����<��"���d��\q�g��,���<�$saKqs�Y�A�BΟ.�d&���{�d?&�J!k��,zL�1�\�a2�i�J#h����N�ua�m��=�Q�ٽ��r�7�Rp��A��>M���Q[���ݖ���_f*�t�S1-{�L�!i+��}V���
�i��1WO�Xw��&3I�\���1����.�ud3�uo���/�m����P4DW����XK��4ԫ��#�c�<�)N1�R�.����O��%<O�we��Rf9'"���0`)r:\�L�L2A���U7К��eG��
�暽�r᠝2qN���ɱ�������EL���x@5-[�ɯ,b����|r��7y���t�a ��}1������9f�3�s� �O���1i��Ǐ�\g�RB�E""��L.f�,Eke���=�#d2�Ho�鞛]�%_ �AJ�gˁR��"�R��ĸT�+�h�Pw<�2fyёd�Q�3���9�x~*�|
q���!S�n��CrsI���|?j��s��-,}��H#�Ф����� �>5���Q�B������wY�D�E��1j��wf�OD�bXs�*q僢6:R��E�W��4ʤ����g�L)>�V��ZG�QD��
�"A+����U[R�Mބ89����VV�q�B�v��J�SD߇���ŮO��6
�P�6;ʛ\q�<��t	q� � ǩ k��^Z����Ŗ6Ag&[{m�b�^8)���b��$b��sj)<qV)ȣb}�)��g��ٮ�B3�I��q� 㒺|����Q��:���2��L�,ۇꯡ$���c]MH]�rۨ�~0�J0S�J�����E�>�����1��j("�;b	W��s�{8+4���2EU���U���"@�}8���G�cǬu�*�E�-����e�N���>����/���<��g���PL鄩^�̳�o�dTXb��"\P��A�+��5˅�m�{ЍSqL4.X����� �PLq�Dȁ~��(�V.D�8����4�dr�\9��k6E:��I��$����3:Y:�ku�1G�QܱP�ѕѼ߯�JL�=X<d�;�1oymO$�g�Fpò"��g��$�6R�cx2z��M�)��@�&�Ϸ?@�k+D���5J�X� ,��Enp�	���B��R4E���Gt����58��XC��:Ǵ�X'���%y�8���ܱ�<U��Z��#:�}����犕��쿂1v��Ek�i�$n�D�D�p޿�&g�n���~��Jr��^���:z%A]�G�� � V(���K[H|Ur/7�<ѫ
'[��R�^0+�8p��#I�5/J"[�D^��p�]1$e�3F\����(8I�?�\�TL["��Έ�X������e�6�]�OR2p���P�:{[��}=1�U�g�`wWT=/��*"l�CQ�#q4Ct�Kh<��h�Šj	Y�ϗL���3��tp1�Ef�Cl��ܫ;䱪���ci,z���q��<YߡJ�/�m���|"Ǔb�%UM][��Ӎ#h�J�Y�)�V��:�7-�QKq�J���yb�qs�R��M���GY�ٔ��c�1Mn�G�K��s�:A�˩Nv�ɹp��i'�-�g�K1n�5�t8�w<� U��[��c8�W@J��Mм�v�SH���j�yi���\�E%9��$���Y)�O����)�2JP��y�_WN)�+.jq��Q+�a���HH<Jlڎ� ��ߦ�ټz��"f"-sm}֭,O�yΜ'F�u�rNF�Gs�Sn�#c}��ջv�N��bAE�"�"�V��wμ\<rh�Ą70�N�4u��+aE��%��<���ǡ�r�t�`�c�q�Ǘ�f��w���1|'���D�S�b�]id6��F�t"n(�#C)��y��� @����pS��G06���Ή���r�RǱ+���*�Is�C�T�O�ҁC�5|良���F�QSq�����Ն�^���S4�t4��*�	���s����Y�D���W-�w-&o���-6ƊZMkl�����|��hV�~<�C�M�M����M�N��U�&��QtȜ'Z<4�� Ԩgt��ꍕ"��^T��Z:y�-�6�q� �k�S�Җ��/�?+�v�����c�+��p��
X�9�#ӛ�$�g���Z��>v��p��L�s�T�(���o;'*H��4�nB_$���vx̤��(3��C�|M<�8���]+K�v�]by	lDFe�S�~�x弿Wt����;�MX�d�KZw|��e�'�C�&$0��<�7D𞨋 �E�(df��v�5.Ff]d9�P���1������Ds���C��&r)����V8 r6���WWW�b��Q��("��N|���V��B�3�!aE���	���(���(?�A�p�T�X����A @�p��*V�9�D9�9v����0.��shg=�΁r�� ��"�����NiN�3P<2�8��F��GM�!#r��I稩�2w���[oI "��=s��t��c���\���}'R�3�$Rw�����m�=�L�{#�#gcl��ɋ�1ǌ�K�\�&�$��r�5�?{¹9Q�CU�ND�"����8�$��㤽X���}W�s�5Ǝ����8�t��\%��;oS�P��ꓙ&��t�Cd�W�CI3�������&',+uV)��ȭܧ�;�,�$�ވ���c������6#�3M"�'|�ͪBQD�S,1Q�S&wV�Oq�Di/+�9bI��Z^�Sg� �g�jWT�F��)�B�K�T��y�������CD�sD����S!:���/�]����䲑2y��L'j0��r���L��sH��5a=���F��R�e���
*>�q!RS��/#���\�8A���f� �d.1y���u
��{Z��@�&Q
����?���1���*��v6|�)�c��9&9."���=�\��B�k]N���:?C��U_� �+�l���I��r�B���6��f��=��1��+��@�CS�������K\�Y]�E('�ͭS�[�S��Nl�8�H��!��g)T��4��A6�r^�M��8�U>g�a��T�;�˼�C4LΣ���.�r��Tnju�u^Vb��4ƨV��.�A���d�$8�x:-ST͹�N����bל$����b����F7�cE��|�Ikݼ�����&��B�l��+�^��L���$ }�T�л��^���:���"�吺ʔ���R������F�)�8c:,�צ3��I.��M"Ӧ�>':���&��?8�^���cҮ�Xu(�ܱ��@����M��Kk<��&�����2g��U���c8�\A_�B�gd7�r�/�|U�J`�j��r�CYk�:SN@��e���#��*���?a�uF�p>�r��Nv�N�2B<�Ek�J��f{��}*�J.!�Ѽe:�ܦ��2������S%�9�'�E/|Py�cps�|S@�g��	gb�WnL�e�0I��Q��4�i}����;t`��ϝF��Dz'�s*�8Y�WS,Ѭ���p�J�kEC�q3anɤ^CNbZN8�}����309����>�:��aV̳-f�f�	uE���I��.��gPQ5Itq�YGIg��M\�$��A$ЙM�M�_uu?/�6x]�+"f �5ӵ���Q�p�W���!�7��ʞDD�q�%	��8�p����� f�1%�2�43�D@.Qi�}Nu��NG9��Fky&�wv;��J�ce�i��ƴ��P~C-3�d��Y�}b'����l�>17�M�>��P-*/�}���Y��X*	U�C�a�+�G�cU���4���ݦ0��!lTv���(���'�K*���=��R>��X6���袧�T[*��Y���)3A�X��)\1d?,�a��^��,�w���0��^'���E{�#n�ZAE+�����>�vJ8�����z�7WP&S�Ӿ��R<��R_��Ϥk��<��&�TYt�Y��e���z�}�F���ey���	���5ϫ�`}��7=dL��P֩�t'2�P���0}��44ϫ��01c�1񙓝;mY'T�odx͋<�֐���)E�	^��!�v�~�e4�xf����i'nSI���!L�qvR���ʛټ��:�d�g6�}&����x/�"�N2����X��
u�N3�b�ݎ��fI�;nF��+����Dj�Y�S�c+}(W��c�Z�����,�3�����}�U���ѱ5Ь�e�����5�ډ�2KR
����I��5�:�(���LΒ��o�p0�`��NOXR�B�'�SX�o�4��Q��O��y�:�vS�B 3����ދ?�x޵�De�on�Ç�������O��޹X�>�\G���mNb�'�"�/+�W�עs$�����ZT)�?o��Ҳ�Ԏ�~��w�g�Bl�x��y�o^\��\2O!���_��>��o_Y�����ُ;^�QH���$�s�>�G�I��8�R�~�6B�^���ksp��R�r�%TV�7v�Л��w��%�[76�,�x�|�jg
�;n�܉��է�qY�Ƥ6����m�~��* ���*͔!g1�+O��޳T��
��C�L�#gy�/���ۨ�~�X.|�a�)��������}N�$s����� Mu�y'�h�y�K�:��7.��I12�0�\���o�Kp��K���o�FQVЄ[����_��ԃ821W�f�%��"4�Ǖ(��<�L��܅���Fݟ���n��m����D���W�êP���?~�"l�?��)J�)�8^O1ű'��B��_j힥����e(�ĥ�������W����w��l�,��w/���.�'M�՟��^��:���&���&6���P�߾P%��գ�0M'�����
��=�*�g"H��xa25S|X�I@���RE��3G���U9���mQ|Pg}�6����G��j]���S"2���"�&��Ay��/���:9��Ib&�Q���j22�g�7E�p̔Ɓ;�+uK���E�E��t?։{��s��~r\���M�6��x�[��M6��>�)���1��<�>Ӏn ޻o@�R��EG|�:T�����l[%Y?xpI��E?�j��������{Dq
E$�p�菜I�����JI����|*U�D�l"7�B,�o�������v��J�_�����_�E"�9A*рOOo���VP(��T�g����bi����)*�+b�Q��XS�RN?x^9^hUȾ�*{Y��cD7�N���~,���xE5��X���#��gu)>q_�B�gO����`O���l��c%	cgg����-dr�����d�"�ơ㚊�"�8R�CB���I�)��N����$���[*q��P���*��xn8n�<,CD���W��[�T	�o߿L=����̯����O=� �C��j��G���fU�N��ߥO*�|�Emh3Q9���g���˰�����7ԙ5��
���dm�/k��]W��U9�9_�����F�F�����c׿{�MM���\��nb�g^2��_D!�}��Fu�5,#�=�0g��±�:�~�_	 Y���OE]��ͬS'`���#J�(ȉ�W��LGr�i�K���i�q9	ݓ)c��o��5�
���lD֗oU�3ǭ!a�0ӎ���"ޓ<wR�x�2{�a�����٦���?<ێ��ܲ��W�s{�hVb�xm���i��3�9oOs�#uzf�T��[�55�K۸�6�w�"��$m��xjl2]sj\��M֜=SRx�V����Y4�wwG������h�09&r�L��3��YZY^9W���NS�M2Փ����~�w ��7�(<�&�Қ�\�����@��>�s�)K��[�����3ճ&S��-�p�3J��B�D�h�T�P�y�D�ԍ�v�J$�|a^1���W�+�T�����Ɯ)n�}������39#cR��BF>O���@1!-���֜����[3aA�e�)��_81��Q�b� 3z�hl>�i}p���v:B2ݓY�\�$���`��?��+sN*.a�6��^��8A���`v$�Z.�ᆚNQ,� Yv�=!��gU�T���d0&@3��Y����u���@�b���EB��Y������k6kcXf�d�;,%�X��0`N�C&�q77�2c�Il����l{�)VÊ2Mm��}9xn��F�6�-F��,�c�1�2��B��$h�{�Ddn*L�9U��L��@˄+����\��ؘ��N���f�EW��8N��`:-+"����SK��}Y���49x*y��!p	�P+�R�������csӎ���-�BB92�Y��Nuc����2�c��0�6�����lSz�[�MA�yZ(�cL�Ζ��z�Ck��&�0M�������i�\��������2��\    IEND�B`�PK   *_�X� ��! �3 /   images/646dce44-14bb-4c05-881a-5e107587e346.pngd{eP\A��������݃���u��%�BBܝ �%�Kp�`����߭�����vg��������5�1���@ ����.��!��B�	���TwC/(���.��^�%�����7[o?O����������������	2��� ���a�A1��T=o!�Ŗٖ���A���GT噧cԅr�k��,����vH58Q�ͤq�������Å3x�HI^c�P�~Q{��gxei{�v�Jv�"�����pI��í�m��͔	��8�g� ��v)�Ep+uc�aʪ�b	D���� O��8x��A������#�֟���OQ<#�����F�[�<Q�kU_,j	����},��php��E�l�z���:^)�����z�o�FR"��:���y���B�	��.���'�җ9����l�휗9d	>��z�w�/s��#�Ү?��@��C�]��s9�����D�z>�RF!�Xj��h�G��rѩg[xq�h��2�i�����$id&�`EQ��R,楚�Pĩ�W^ }��ƽ܅c��??���`.q���d���/*�
�9S���L�(���{���8��j��ѹ���b��Mҥ�����U��#I���ջlA���G�,��ϐH)l��̑�������Ļ����Ĳ!��jV�H��`bG�ϻ�2.q�",̮����H���r��1#��OVp5�-A�[��%��q���H��]���<9�6��&EB�(R���n"0��_�մ�9Z	b�@���&�ghk����������.n��x�}Z�V����!���UT8���<<
]�`����s�ǔ���{��x:_�7�K�!���B��Q:9ځ�)��+Gг����蒖t��d�E+�^4j-���?�|b઺=hzQ�w��)!�nա�9��
�-�W�_kVg��Qe��7et�R����edע�g���T��{T�q�O/dՐ>�o����5c�,�����}xW�$x�)o��_���ƈ�8�2�z�#��7~hP��4�h��}�/���'z������و��ޟ^r���}pCY�E��~� �p�J���Q��[�y�f��� q�+FO)#�$���9)�Y�����������o�*�*�����]�{�3���Ji�<�e�y:ɣ{��U4�bf��߮	͛ͮ��e�i�<�#����~g��Ro(�8�EA�{�`��A�������ټ6JńY�-+��+��ȤX��o֚˙���6�J��}�	�`B>B:�_uI*	�����VB_@�q��������r�����l�����7�t�<�D�ë�uD�Hw��jjǢCS����t�H[`}KL�O�38����݇���R@AzE�h�"��n�T��Iy�.���.���^y
?ܲ��f�;�i�3SU�N�Ä��	��{J��� �z�@�������[s}{]�,�i+E`ЙV�:�y����ïH��wy{)N�o;���^<l�~Ic�
�������w�Z=%�^�X	�ů���NWD
�j�d<�N-ۮl�
{E��������|����=���?}�"�$� ��#���(�vG"����
��P��?D�zr ��j���`�����l��0e�z}�~X��q��S�i�Qʸ���A��a%�;>�l�5EG`���ul$��̍#�EOC5�G�>}�Br�0��8�"=L�o�]x'�^���wxz��~�S���.��NA�d���Z�p�~4��Y-Ƕ��=�L��q�̸WO�s�*{���Qf�)%��H�¤��:���� �K25��eË�%y��@q���	K�"�ŗ�c�/���4���oxY�[�	ت���"}?>�eF2��(*8�@&	|���%/��b��$�m�
@V"�83�`Q�������c��D��Fx^,g�WeN�R^M6Ŷl �j&O�DE�^���� ʍ�G����s��Ʋq��r��xVa�*x=�^�pEt}��҂���k�$/�� �K+��v?I��$iߞU�M���2�;�;q�1��b$��a�,��[څ�f[c�Q��Ř�(�c�����ڲw!&/c�3�������Tm�㉗����nW��7����-��r瓚'!�`B���
���>Pb�a!�������M���p���u/pz��Ӵ�s�'L&2�&�R�MY?� ���B�֞>/̂+�]�����`�R<va�LZȟi�*i=���)z����ē1|Y�D�"�QA =�3�`�2�b-�����r�/Y-	G��tk+h����^&Z�b3�I��/�M�@}uf/�ሺ��:�b�Y��x����ǳ��զۭ�^`��<II�L<�ۖ@��z>wD�:I$1((��{������}7�.6鯿��XdYX��J�;���h����0�1LO�78
�����������5u	T-���?�œ���Z����Ya:r%��<��W�S���i��e�0�s9�hi��I�)���OU��t�u���6x���zA���}��l����d	�1��ˀ��7��^����S?�ʺk��O�bG�����3{����⬰�pQ��Z��'�7�s����J���=������m����$�Nrca��Bn����٦4�cЅ�(�nTTACz�� bg�ϠU)�n�2�g�kƹ$��_�ߠM͞��T�u��R}>!�s�U:��9�����y�QQtLEc�wT+,����W��s�7��4v%:#JmiD�ٕr�2��S˲$�U���E����5�C�e+2���B�&��P�?8q�ʘk�`�0m&9����9Ë�Zﬀe'P{Џ>�N~y�aܑ�,���h�>��cY��E-�D�x�'�Нv�O	�T�u-Q ��$�(Q�4-ZI��ړKI�J�ײ��Jr���.j�Z�L�#~%�J�s��&fEyq��yjB��?rO}�i2��������Fz��_o��(ŠId2;�P����q��@�Z2&�ؓj�F�^	s-��u���^ �xG.?��d�5���W��+�|��-�^�%{92'��z���K]V��O{ou1�N� *�,
�0~Ca�(%�?��-fx��*�b�= ��i�<M��Kc�z�J��b�'���Mw�d�3�*@�&G�_��*jW\�:�W�z�"��hF&�--�^�6:p�S������ͫ�N։��KL����L���e�R���2�� �GǸKǵ�^�^ u�H���EJ�#�����V*�	�g�m�����9���"\-���%��d�/���#�F#ˋ[6����t秫�wf�ӮTF�ߟ���+�G����H�`�mW�9�X+:�K�25풮���_���8�a�
&�G0�Ac��.hP5�_X�Y���b��]��0�޳	�K�#a�54K'�
 ǂj-F�}�z�
�totIo�/y����b��5��!�h��T��D�������N�݌�r����ԛYOʸRnIJ�ym�-���g�:�n�I��.WU6E���;m������6����T=Wb1igG�ԍ�~�h�8���}�����D+	�#���Z3	�w͒��U�^Hc ?�jn��p ��|#������% d7$�Ю*ǝ��4\)V?TP��PbW�mN<���'ؑH�ZbջH��,�i�����!�����]���� �c�3*��Z���tG���pؐ33dS��Tу���1��s~�>fd���+�	����_�ӓc��?�.���b��УA��;+�����I���J<��am'La�l��������;���dͶ�!u���
x�]��=sSq�UVi�Qb_�M3��Fv��t�6�J�Fv-���fki�B�('�Y�FJà��s�kiW���P[�p?4		�Y9��.������֙x>>V1�0`���TNLSd��y�0����!��#�v0��E��%<TK��,C��z$�6�}�����V��A
W���y��P���������W�G�2'r������Я!�Xǎb���o�Wﻈ��1FZWi�\�Q��_Κ��JFQ�{�׻�:Q�܋�>�?ny�"*�U��#��?��r�FJ7Q�D6z��5���()��E*��708�J�}?	�`:�O�4�4}��1�� �F����]�@�Lͣ�L��ۊh�����|��F�4��ݥ�����O-����-��誰��!��vOr;͇���1�0�o� -:�l��\d!���+'֗O)���wͰ$�L�S��Z�,��/`���@��{�@@bA���9]��q� ����Bˁ�7UeݭQ�YG���s��=�J������GN�w.�E%/���v��/����hʡ[�"Ek՞����Nt�`�
D�������H!�GO����S�	;�UP��t8b� cL�A�=MG���' ��T��-KH��KG���:)e3Y����������Xw��mĆ�����x~�����<���l����M�}��\�`�i+��M�gzu�]�ՀA<��Ԣ���O��4L��⏢����cɋ��7�$_%���W�
��n~Jh�/:H����|�')7?���'@�|JR侄)L;����R隭�����0�/��n���W�E�ܢ��&�E���{�Oo��|d��MM��'����\���c�H�#�c���?<�2�Ua(���}^��"����>֫�����U�k�nK��l&�K�ۏ�F�2�fc��$Ǿi@}�c܇��.��)��I᥃��И�a�s�-������ƿ0���9��ó��_7e �rſ���!����U� Ds0E��X)e��i���-�8�b��O�؅~�1"Be%ݼlD�\^��|�4��E#���є��uV��"f�_da>���3�!�8������|D��_;l�"Ҟ|�>{z��m����I���i#�(Mx=�5��рA�Dq��?����7�y~.��C�����!�j�q=]O~��^�}��-�L��eaI ��.����{��sH}aB~"�r(t��=fW��u}�z�{f����t�΀F��r�ZHWtB>s�i��#�b~�L,z3ܶ�|31Y'�x�k�:m͕Niɩ��)�f������O�3��o���I�"T[�J$���~U�oh�B\�Vx���X�����LK�����T���'���V�o]���܂�ECM0-zS�d��EM��c��â��n�U�A���]�J�w�sg�C�}��P$l��:�n������U^Z��P���&���o�-��w�6���W�Y�Z����|�jU<W�|r��:,�B8!vcբ�v�#�		�d�a���)pۢ��񟔡�_1B�&~���e�shF��.�®+��!|B�y������R����/4�L~Ws�fЅY=��3x�/��t������߇@_��kv���{�����@X�˟|���H��1����
w��#��ݼ1f���Đ�dv|i��47%x�������A���a�=�K�E��\���Y�?�m»��A��ju��Y�eD�vE�~���&�1�ްXڏ{�s�tD�y�ῗu�mK-z��廪��ɛ���L���2�fd���Zb=3^J�!����Lzc����#���	C@�B:��η�Z#q6�T\Z����M�f�Z��υ��nd#YX�$�󀾣��V1Moa�<PB.o��^����%T^�ڣ�JVSmC��P4�*��󒿌�^9A��Jbw^�6�滚����]��M������4��A��S�y�)��.�����j�+֌�2M��*L���X��_K�|&;�^V<��,�~cͻ^�}�߇����53��P�ճ�Ɩ�E;�8����Sr�KJX�\����.-g����i�4��Tp�"��@�M��)K��mR��(���I�>��]ރ7��?z�>8T��a�N}~���HU�Jh�WX�a��LV�C�-Q+&w���x\����[��b���=|nu[IFӒ�����g�q|/�n��G�^�	X<|�b��o�w��n�'��8llC�h�����I�� #�Q���`�����Ev�y�̫�=��v~uRBu�-\z�$�zf'!�ی�KP?rZ�J�앯�w���k����yH��'��K��Eќ�G�H����@'��#&�����'�R�.��Lb��(1���)79�aq�!d���`!�m��<��S�ו5�dO-�E��\��P��4:��O~e��^�͏�Z����x�pW�]��p���B	������-�%V�*�z���w�����iiy��{�Q�'�c'*���W`2F~�w�]s��`��? ��8��+���#����~GԷ�L����fm�ݝ�e���C�[��4�_�����0/�Fxu�<j�������Tw�Rf^��i`4f$ ʎ)��px�CNW�)�'����"6� Y�� �P~�,�,����Ik|���I�0]�5 ��҈��t�d�d��m���<�q���C9�k&���;v��K
�Di��	o��Ĕ�;"t�̥��߆��`D6�GB�R��g#?���0-���%M���c����8N�+I���FH�8��M���QGr��1�9���M&4�|��<1\Ƴ��S?};�(T�QRմ��������Kj�<UT��w.9��Ƃ��W]|s���մ�`�ѣ�ܨ��IB�}o9��}+wa ���)A&e"��S�f]^}ɸ�'�i����kw��4��Sek�L\�_1W6t�Bo��_E�X���~'����=���>d��$�C����т��uj?�KOԬw��Q=�I�H�)����4��k�Snc?����0W:)D�Us����.���T���L�Ј��א_�`�x�9U��*��?ކ�n'xe.�H��IbG�bV�Y��bw%2�`ǝ1�F�ڷ�����QKV�
{xd���ț���Z�<���\5�����oY�\RWry���J�UT �5���X�EE�	�ӫ ��C��d�� v�?�k�%T�bu�����ܪ�� ��*E�4��ߑ�]�dIPۥ_N��X�񸓼�n8��6��7�K�j[�G�B�]T�W��N:�}�[�*�1�;����Y3�;��.�Ru뀟�"��~-3:�ug<��g�L�#�I������r�C��"�<�z'��뙼�ET�(g�hP;\�8�q�͵��9 �%!�Y�O�����W�I�0+�"C�v���]�K[KLܽY�h	ie� ejf�He��������[�C��]E�� �99�>#ۍ\���tq��fW�#�������p;�[?蟓XmA;F����awjM��w�A���+t��!���Y���nץnt�!�1�b7U��c��.��<պy6�)��3�giQ
���T���+��k���J�v� ��[���Iǌ���!�N{���zQV��%L��^������@�t����|1��� ~a�}u�)��1nt=��2�#��N���6�9������Q�IDK��\��������Pǭt�η��}��v$�_�[^v�bFKk�Ƹ($���ͧ��e�'�6�x_��9�F�ږ���,/IBI;�lQB�N>@�U�ȟn�i	il�mOL���#u.��[�^����:��$!���^�q�䭭Er@U�P�+fʡ�/��Ao5Y���	2�����p�Y8
c�#ؼ}�h֙�bH&�p��ޢ-���O-Ufs�G���-{�8�M���c}"T�d���} 6V���M��u��H���Y�=13~�����*�Qyu�v.���Կˋ���T����D�����C�ώ��ꂴR���>���c��]7/�e��9��L�g�
Z��1�h$�q���V}1�60f���I�ۃ�=37}����E�vtT�W��Lj[�HY6��f�cG��f��=x$H�La��ub����.���y�FLR�|�N-=��v��_T~?q'��9GnJT�޲}��D$��m�rb������v3149�(w��ܩiyV������Y��P���)��RĮ��*V��[��_7i���8E揷�ڦ��$���(�@{l�"Z�]�#_'9�lO�o�cж�T������gs�)�LH<ұ�����g�����"X�,��Z���E������|��ղK��0�}	�17^�z���mVq�!��?]��W��2�rhT��Ր#�`W6��TX�Ҧ��mZ��ƅ���cn��Վ�<��O���r�|-��,[�,
6Hˠ
�#�|HN�w��W����(>�-H��{��c�%L~(�+��J+��r��96+(�	���hל6ͪp�H�{��{�8��E��B\_(����t�*{n�6�ݫ���
91˵7�Z���E�6����ܦ�?g��՞��j���PY]�~��_@��囬���̒�<M�{D5��{����J���[� �!��7��񛔏�c�ba��}N�)�����j�G鶬�1S�٬L�a�%Ҙ�Ť����\)@����4��������lV؍��m� �E�"9/�K��b�eC��K�qw�t��}$�W����g��{�����;����x_��'kf}�u��e����1�U�篆�k�7�|<�+j</�I)����P>d\�����	����ڧ4Eq�xvW���l�t(�z�:�H��=j����Nf̉��F�F��͇��o�!C��q�" �'�����4�5�[S����w+)�=o�ܔZ;
�9�Y�Q���G3����W��a�PV�	�@%�z- ����&¾�gb���*g�i�'���$#�i����_�J�|�u�;��r;�T��G�q�u!p[���v0���ܴo�%5�8P�L! f�k��z)|���o4c��c?YP
^����M�EHg7�o�07y_���2Ƕ��Lj�w�S��m�0�_�Xk��DǴ+��v�
���m�KO�<S����U�_�o�3i�FP2eO"\絴Ay���0���4�86y��QW3	���J�s�zY�����8*TX�������0=MG����(��(#R�q����a,���(��۞�}�0��6�wC�ߖ��0�F[���(��ٹ����b�'���j�[�y��k>���Q5��mqVE)��:!sC�[�3ʸ�_�4u��K������(�C���`j�V�
�����J�4�������<~�O뾋�cl�v�Xt�N���~Rn?���`�
�RjHV%Mu�+"�2�����d�K�r�eF�)A����nL�5d6��q���m��ʿ`:����N�g@Q�nqF��J��}2,�-p���F�.�t����^�@B�����A3(�������j�6���@��v��#�Ƚ1�T��P�J�q�a�	Rh@�k!��mNR��*�V���Ns#�;5T�K��Fd����b`>]٨(��5��T�*����;���Դ��.�V������:����#����vO�1C�M͗���1�%R_�O"q��;(G�J�5���c�y�1
"�ԑ�K3���]"�F��1��gM�f����E����[^[������xݾ�z]4�n��������enNB�>'!���KԢ3��n�5v��#~�L��aJ��������R���5�[�^��Ư#yJ%փ��[���=[9
��;�i&���赏(��>p��,�]vV(����DV�kC_w]&�!��.p�8��8`��-Q��vũA<⢨Ǻ����o�m����=�?�~f��2o�+Ĳ5�ب>��`*K��~��X���m;�ʷ��n��Ն�6w̩���a���&e(�~��s���KWf��0��ϧ�RK&�2�i!�zڊ�ay�H���\�R5k�Tc���Ц^	",�,�h<�0�7�����}�~/���Z��H&)��5�IY�
��� �hDY�F�E� ��;�m��`1��⌳%�i���o4}x~�Ti�2.�)D/�]�U"��(8 -�}�\5v���i������:�80�,Z����	�+oXJ�Rs'$�;$?BE�i��y\�ZL���ۿ�������sn%9>�^����p���kt�����M��'�₳���T:�~R�Jz`'$ŏ/����S�	�9���=�{*a��+Sd2���S�Bbmc�q�	�/���*����k�x5��%_V�>Ӱ/-�n��#�ɠ�R�W�6�����23�9�l���N�e}x���E�˱\�,��K]����YG!Ʀ��آ
S�xu�H�-Ȫ*�!7�L�����^��
��xS���PEl�Di�
�L$v�N@���592���$%EKEIדi nxC�pϯG�~U0�)�"�me뫪���T�2=F^|������Pl�������)$�^�!68XL���!]���N}\�j����"���0qb��T��K";�?�����E��Q�l��DĲ'�pމ���v�*zH�n�R8k���n.e����%3O�(��]�K$�8���`���@��X�嘯���=v(�44��3�<�q6��?���]�:�M�����#�(�_q��0"�p\����+Q׷h)�"�
Jf�Dr�B���J�Q����x]2U�zUO5��s�
���v�̣6��m��5%>�BA�m�ه0�*�pe��e4-Ҥ���RW�U?�DN�F*:U$󎜠��(�?aj/rG��dۊ���)�Ψ,w'D��;��Kga�i_/K'Vx�A̪R�����9��J8���Cj�]�^����|q|�����N��5�}�&@/�M�"M�>Y���]�Z�
�V�ZU�A��u䔖w$�$sS虳'�/C@�s-�ȣ0p�Ԋ�H�6�q��ǩI 6���QW���"�	r;�}�9�ϰ����(V[�YG�RZ�K|���%~?Ib����@�*M���㊭�3�iz�]"��:V�q\J�����al�t:|>�8��V��A�u��<�$�q����@ۺ�
��9����ީڈ֐��OQ�~&����?!Kۛ�0zg�)�n����`�Oa��
��n�O��}��B�?6c��G�8���1�}@������!�9E�e����|�4
$ݲY��j�D��I��@��K:ڱ��0�5?F�}|�����#�k�a �p��x�;d�z�<Qf�O;J�| Qj�
n�=�kOj��.���[8Yr���(��3��&L��Я�_�_t���T��L>�rR��'���ӫ�몢�4`>Ja/�GuI�A����B�S��!
��!2wK��%�,!q�ag�)e.������׆@�}չ�T�nY�a����7��oUVGl�ӱr>^�T:���O��8=/� �78�{׏P���:�^i�K��u�`޼�*[�*�����t6x��d��\�WQ��0��x4TB�C�P��[*�Ph0�_���o�g�@4NE��*�:!��6�=pVLp;�����i#9�!RB���!�a�lx�g��Hf���J¹�8����L�e�ƨ���i�D�$��gQ��r� b/\�8b�-��)�.�!Yޑb�~�Do����3��?�Qhّ� �' �a�t$l-���-��HB�R��T��*'�p,�^�]��Θt:��-B�rroMd���s�rãx'�~F���`�S�"��͠���)#L�?%�!��E�E��Y@�)�<��m�-:���>E�z���̩�N#���A�ސ\X�-�KBTga#$���V�����f3���Sd64}�v�k
�29�QSҢi��e�:z��B惛���ՔOi��

Csl��9XI\-��̧N���e��1�-�oZ����A�Td���7�+��0zYn�/c���&�48g%M�X����jԄ���=ƱR��d���ypS��zHd���+r��Ƒ�̏��|fƍ}�du�~}c���&q�sZO���G���7
���S#t'�:�ہ<ǡ���-�f����8�!�	x�\H�<��0U$Y[���8�k&��z����գnY��R��n�f�Kjv��wh����b���֏����(��/0[PB�)���%>��i|j��BJ�k�sM͹���v����Nj�s�/��68�b��*ѱ�!L���Bt�}iZ��n���J�W����v�|��㏁���K�"E�M�LT�5**��������]����;<yVC�!�����7�;�@&'�v��s �U�7���9�EI'Vj
+!HUYZ_�$���/��:��`���[�~�MU��U��K���f�e��vO�!S��/�N��6܋s2���X�z�:���͚��3e�':�2)��My�y�<31�� x�N��g>�5�5�v&��_c���0n����4���4?i��L�L@��\���	`O+̙��H����B� !��m2ݱ߈Ǧx]��X�Ô��QA8Xd�d��g��w#���޾(Z�IP'��ܕ�Y��՞cv
�A�yq\���
� �wb��=�L�I��y� ֩��e�� ����
A�3r���"��S��j���
�����W�9%B���^Y�鵏�Sq�HHO�����Zx�Z��C��I���D �͈E_l�S=�=Sx�>cp��|�h�®�D[�=9!K8]Y�F�� I�-M����\u��8�h�wЯ��B�|���ɭ���D�ˉ@ 
�3f�����1(mO@�ĥ�����ئ��@q0����E`1���T���L��qK��`\��/}���^n�` ���i��8BO�9��Ht���m��%^�^ݍ���j,"�	�+�C1�� ��~4���J����D��Rrʋ�{XM8(�f��|W��X<�ߎ�N�J>��R^"d�rn�n��;3��(ʞ�Cy�K2�Z7�I ���#�c�L�g`��#�kݽ}�`o����#�G\)Ξ���"�������'� �j�G���S�_P�#����.q<Z���џ�Z���dȰ9�	��n.�k��w�%�sYn�~�-Xrs��j�M����e��A&�Q��1f�M?�=�J�� p)��9���IV(�b�J/?�mŮ�J�6�iҒY�g^��	�/:z�;{g�74���æ�q��ӼtY��4��hϭaI�1��řD;w����?��a,۷�V�,�ݞ:�;�q4�T/}�X���Q�+`?�QgdoJ ����_�Y��>/স�Ce��iդ�����0��n΍i���ز��m�*�UQ����q('[����|Ӄ�f��L>��]�J,��3I���S��fN4�Q�<M�A��[���V�����L^|��� M~-˩b�6�`�ɾk��R
9VE����a�9�,s:���H29ֶvP���0>���ۮ+�s���;�ͳ��]�Ԋx6�<_Ƥf�
���-��eu֊%������?�A\j۷_��K���D2��W��.�5a��%EII�]���	�u��l����xO�{�|�KM���ۤ��A�>V����h؄Գ��Q�r��uq���`�n����]�g���_G����������<5��ޑ3	�(��o��G���(�uS9� �����v���iY.f�C�Z��z��h�=��4�/!|$Y|�\1�l_�+!��I�lp���]j� U,���E<z��y�P���}c_��Xo��"��R��"Ķ~���,}�J�ː�k�nl��f	7����-E6mN)P������$ F�(L*v�T���w���0g�[/��U�E��h\�y؟R�Ս*w�T��������};+zF��<���JBMޛ|S;5���f򥟈CFnCH�)8؋	\��&X8k� Bk���l�ec5�{�r���{Qek�hf��-!҃t %1,9/�ڈ�{}�6T�!I���JxY�C�����>�����ֱ�sts�遌
�H�c�5���I6�c���G*t�lRՀ����q1�d��*�:���ⱈwG�2�ȯ��D&��Bs��Ӷ� @��E�����\�?�F��w���qNN�R��>��F5ل��<�|8�Ve�fHK�1�:Ǵ�X��"j��y�����B�k��&���_�(�xAE�,��NC�䞫02��|w3�;�Zg"�Ժ��kQ� 8���xA���J��=�O���Ob�zst�2���4<�ӧ�v�VH��3E듫¸���&����=���[S���f��an�-��We"|0�6S��'k��oJ!}E�I�$3w/�Ŵ���t�a�;U�?��Y/c"���4�N��op[��~^�s[�����n�8D�)�mNߍ)�9:X��Y�Q0kC9[MT��f�*���;�joUTQ����W�X���8p��'0�$˫%�d	R_��<��6��c��\)�l�I3gn�(tf��!
��j�jI��(�~��4���]����S�)�"WZak�a�|�����Uv���'������c�(�CKNP�/�[�;��ə�5�@i�Y��'�F�{]�7Y���l��������\I����!�N�L(��̥l!ϫZ�W���;�@K#L����7]k\�2Q��$�y��sZ �ȅ��Ϲೃ�Kk������ҊSk���c*qa�U�j9n��ϖ��=P�u��b~5�[�@+X��|�|ۡm� qx�r�e;�<��������o	�+�:1Ӽ�ӝ��MS`]ڹ|�u��FB��+��)���7�C)�����q�K͵17?��X�I����[����䭣���]L��k+��M�'Hf��"���Yq���Y��/�6q.�����E�*;K�LJ���߸�x�o��u[8���<X�*{��H��J�.����=wq�7Ҫm���h�Q�(`���k�@n��i{5�n\����[�Kfa7lg� �MVU�L�ʺP#ޫ~xz����e:�����)��w�f�Xd�{�֍C�߆6��i9�-I�te�fl��� ���0��G1����A�L��H~�0�V7��޽a��G�s�Z?��Js�	�i:0�&\�{�~s�i���d'���ī�m���?�2�8���K����O,B����q�)K�|�Dv����Vsd�w�"���]�u�26u$iO�,�y*p����n�݈�b/���p�ݛ��µҎ5�Q�d��V4��D���b;�9�E��痤נM|]9@:V�E>��S,>�x�	��&]���C��8�dǑ���|P��`+?@�1��S�Ԑ���`۳�6��/�����wQ�5B�p�-T�q�;â��d����yս؂Ui$�)V(1A}4=����.�,{���t�ƭ����%�Н��g	~�L��	��+�^�9�ןo.p1��@C�*�b$��ς��B;�ՙt��7�G�G�ϭb���/����3����z���@�&��\���"��"/`*Q��Dy�]�艐�·�M-u.c1���ԁY���v��P��0��	�ID�j��SD���	��zy����
JY�!�v�#$��֝;�5�Gb�~V�{�����,�{w�s�].��>M}�e|]I�h�\���i��9{ ����-���!S�g����'}Er@�^��*6௯)� �vO�/��S��S����d,s�bt �&yc�hH&$�h�,��t�=���R�y{���f%�m�fh����=k�z�wH�W�F�@�w�,����/J]0�۩��GP���*,R�Ϗ�G��I�����9�`,��Ѓ��E��Ϥĳy�gn�؏���+³{��T��޹#b?�� K1Ж��.!����|7Ϙ598�[r9�yU�꺁�џ�54�L���݇u�I۱�<	n�6DR$5X=.�>��� �4�Au��懎|��V�+.�s��6t�D��,�p�@��C2�bj�C@��(����`����y Y1���eim_g&&0��w*V鞐�?���_Y��QsZ6��|�T��u��_3�_�K]x�G$�g6�8g��몎ݯ�#�J|�.̯�Ԕ�&������X��cn�'[�G��J�N���J[6���_�$Lo�>1�J�;���[�/�$��ZL5��
�O�,��RP�+�s��y���y���9z�lVr�G)O�T;�B��%BOM"O�n���N6V㈮��d��&�k[b`d�����ǳ�v��B��Y[��5՟Ȑ�ˉR�2�E��U}d��	�8@	i����2��B�N[I���=a���$���S���.�W_������b��jֈsb�]_]����f�s�Ur�dr=����³S�k`D�\~B���Y	����Hǜ	ъ���aL�s���#-褕�k��%H�Խ&%��I���#�K�
U;t��Ŝu��*5�<N��r+D$C=�������y���z?�#dP)Μq�K���J�8��n��ə�N�4�������5�5Ì䉏 8ž���n�o���ܕ�	6R���� ����~|	��C)š:~�����5��Uۭ&QqZ}���8#k�;0�H��������C*�ﲾ�CfQ�vkC����"�gY�����[�E���CI�� "  �4�"��"��(% !�]R���H�8�H=�5���;�}�s}����y��b��^�Y�z���g��'���0��f���:w�tg$�	fV��?8�q^p�/^�f�ym�!����/K�h����-�*���^]�l�q>�Rܲ�����a�I�¡|dKT����������)GQ�'Z�X�
�aY5��Y���QV(}˝�{�5)#�	���k����E������O΅ì,V��F���	[^<�[=͒a��ǜ�x}�O>��̞���}�y+���_i���� xI�8�Of^�=��R�#����ƛ��G�9dD�7`��z�4��8�3P�!�Nxވ��/R�>S����+$�� �.ġo?<�W%	ݘ؝�~|�q~*f������p�Ʊ�Js�M�s�4��W��\�+7B��xc��婙���3J1�����=ϩ<��͍��,�!
M)�'-���}���zu�9�?*�q�x_��D�.�R�A.-7�$��F�]�CU�� ��j�&B�C�ӓ@0J7P�=�+y�M�����I�گ��>5������sx���������;տ\-�"@�k]&�^���!W��Aa]��F*�]O��T�����:�����ٓ�����k��4�}�
�r�r�zT�G��/�d�����WO�i���~��|�<�v�l�?�-����w+�i�]�=^�Y�Ԕ؂`��_��_�<�<���Kq�����>�dm���h�C!�u��/6���gM�Y������`��������}�*G�.�|��~&��u?�MG�R�����J��#x�z��+kF���k(E��<o���_�:��x�智�e��ҋ�����������i�N��g��.�p4|����g�C8y��m��k\��oK���wAB�<�Ql���׻h�3
�����f�3I\�����DLǌc&���:�>7i����	�O>�i��9q�A��Z��m�j��ǴRѶ�$M�>��7�'\�V�4sW�-��!.Fx�.B3g/���~��d��[��!���9�cZE��:RC��8�o?~ӽ�����s��g8��C�[�2�4V'����u�i��.�\)��L7;±!3J�>�jU&��^��=$i��Lw5�_��;����qr��s#u��]�m���"��U����^�_�mb.P����������+Gh�;�%�L���Iy�^Ȉ�v�<�Bh����~����諴\�y���܇��a(*nrc"i+���2N����mځ�	��;���q��^�i5G	ߖ����i�A0����1�������;�>�^^<���G��x�
6kZn6����E�}^����H�P�>r�@f�
;D�gԕ�9�>�dL��#Q�xN���h���W�%e2[�'�>,�g,��
J;�ӘG��?}r�N��0�AR@�Pa"����)�)���/�*ve�P���2w]�>ؙ���]4�M�}y��?�e�W��{���$�9^�8+P58Ny�>��8�j�t������s��JR��I[�����E�w�^��DA�`�v��p��Nwb2��P�����?I��=�ťxwf�}����eTA^�T�7������q���33����x�Y2�� +��-V�aՇ$_p~*5�e���uw4p~~�_v� 3d��B�pPk�%�\��T�<����yL�0�J���]�L,��zDH�ʚN�`�'�G�Jc���IF��3���x2�+�l�`#�~P����U�E�'_OeT��O��A��ʬ@1����A~�'�I�f
!�n!Wt:w�c�|7��3�!�+
�z(sRH��sS�>~Od����x��d�����su����\�/��f,)�ψŉ�H�*��o�u2l����������Ē����u�x�9xe^_Z�W<#�S>�{�G�7`�_f3��ə1�+_��b�]�7������~��L����`�9��[x��Fő`���ٸ�I"W�p!�gx�Q��=�Bd�~�퍻����|�t�,��G��fV:+��*}�U�=?�!�<�	l՛����BaQ���H�Wrи�bd�<e��ٰ�>d�Pr�q���}JdΣ�w���D��C�q������z�~������.?�x�<U��[�W3|6W�RCX>+8�I�ֳ���b��Bw�^�$�Ѯ�t���7yQ����������*��1�5x72
����v��w��;SN3����}R�*]�Е�ӳ���+z2g����E������׫(�`�kg���+�"���0u��%ٺ�u[Qˡ��ʳ0*���j���_�A��'�|_�~�1x�Z����R���U��|`��>u�Z8J2�񙸛U�/��^��ޝw�<kmN{�!����òؑ�<X/.�����,'+�B�P6�佺ƈ�������sm�@~5LL�ި���/>�5�	����a�Z�Ltlg����"����k�5*�R!�����*oK)a��(��ߨ8��F�����7{;ڽ��s��I��m�֚�XݹO�uwv���~N(hμ>k��+5d�[�͋��,˫�����!Z�f�RK�����H��J�ӣqVvȗ|��ɦ���Y
���1��yʭ����hH_�>V[�<P7���a1��a�����.wIN�����'e�T�N1"�<�&�Gz�Zc�=��6��Rm�N~��,-}t�M�ҙSt|].�5������=�I�7�!��:;;nWD6b��n��gh�c��3����3�W��lCms{!r7�Y)Ũ��mZ��n�d:�������a���Y��>��풹�ϪvQ~zaG��^�!qe�[���O�uy?�2�� �?�8tx�E�+��xK� ;)q޻��GhgX�ͫ���0��~��f>�WT���s��	z/,���[�߳}�v]���X�̟�0p�ZW񁏦Mχ�Q��}�n�B���|��K�f@|��L^.�zά��Ҭs���*������yO����02��%�$R&F���
}*���F�q��2���lr/.T�;y ���:�Q͗�϶|��R��xRn?749_��+;�Rϒ��A=��1w���.����)4،���8��fC��r.�uи��$JX-"��oKY�mn���{�=��A�qͅn��"ԙ��l��*i��:��D�4������Q�5ߍi������n���h[�@��O��Δ}wĖm�`_m��f����V`h�������C�����w8�n|̽J���.6-����y?L�8�m�?3e�9g�H>u��|�H���R�~�{���4��18p��dC����V(,��-32�xZ���p����o�2���IB�I���庂�+�:�4�OPO�
�Ŕ&�>pV���*�L�FyZ-g�Vg���F4�"uTD��觳���ԥ^i��M1��<�d�,u$o�g����Gh�_ ��7ܭ���Y��8�0Ezܾ8o��)���b�W��}�k�j{�L����H��ݨ�{�Q�kˇąuII���
���[���Wδ�5B���G)V
���O�fs� �2��[���m�@<����u�DK.Y�����&j�s��=��d(.�/�yA��.��V�X�Ϙ����+j��]vv~UȜϫ�0�D�{����p�������
*�=,F
�'p�X�I7�9�A��^�R�P��y�f��vך��Tp�u:�Ή'=]s	�T�Uߢך~]1�F��5�Ԛ�tC��l��/�߄�+FL��~Մ&�3�3�IM�y�*��V<�[J�$Pa�Í2MW��j�����Q®=��R�	��1��_Y&";T*ag���Ψ�4����㠒�eq��?E�V
憝&�%�x���Jx�,��"gv>��-�=>��[M�zHw(�V�\8��q�ҽp� �i2�����.U��<i�%7� �y����=GM��3�.��MA6�F���H1u�b�z��W��a��r�FT��9s�w��z�X9�A��������j`f��M�؈��
SuY���l��!�܆V��wLl�2ڙ�c6ɓ�9�̹�6@��*�L���Βk�z�=��:���n\��a�<٭:*]�<�G�[0�*����S�R'�:�^�����2��㊾�����l5�/��N�y�X�.�0�v��x��=���V֣��zkL��=��ъ:�W����D�&�S,��4Do��Fz��n�r�	�ӡ^�ae�63��qyH+�~�$!��9��j2&|��-%�x�So��J���v��,���*��s�� ��T��w�)>Յ�9��#:��a�fS�j���:�S����7ɎH�ڡun{�����R��`��7<��d�R^u�����9����~��P��\NY���M<,��l �%4�#1�5���L�=��>,�T��+�[݆���<�{(&�^.=�+1����s�ݨ�*)���;ߚ��T���q�R��!c�rI���I�<ϟo߈-
��,��	��"v��j
!u���!��n&��<��/�W��>�څ�PK(yY?�p�v98K��s:��Tc0vI� �(�0�ô���o�P������m�+����/5�Ա�>c�^���������&������\o���d�|kQ^d.Z�X����}�u!�2�؀�,��܉�Z ��V��=�/R|��F��hc��R��d��Ѭ��Ng�!�Jj3��[�%vp�Q7\�A1��9�������W�K����f�uF%e�.*�$�����I�\*)Yeٔh.7K���(dGM�ΜK��)�\K;�â�0��ץ�e\��Y�xK�]���;�e���q����%�x4Vm F��n����/��$T�w/��1����r� ��"*��i�\*���#3��)�^8�J�F������G�_�l�:%��hE� ��&R
ȥ��~Z�P���f�Y��S�%גU*#ZW�9]T*�5m
c�����2����˖�Gvg�y+adL�e׏��T��2"��g�$J�~���1<�q���A1]Dep�j��"L�J����}�t&6�Z�<�}���H��.��~�n���#�;�eP�����+�u��#p�&����3�_���r�}�M1E���6"����c����Dy���YX��2�G�W����R�(/�?���0��j��Fwp��.�����n�������ƈ]�('��8޶%�h,��$�>�a1�c���E�_�-H�/T�,��Z�Zp7�.��nPW�BZȐ}��Sp��]g�h���1f�lCm���ѯ�<����Z���!��3JGz�Z.g�D6IX��o/��/��kf.���^�q�C���g�E�%u�g��);eNx�>�E�̠�������[��$8����!fĪ�l�u�zDt���VMqbYX(Z���Ä ?�%�r��}��CT
��Ɣ_Pv-O���|�i;5��პ��:ūJ������r_o��-;���.�؏�h_��xI�c ��ٚ�;_[�<��b��ݲ�"VyCz��5ake|~����p0{�O;��&�(/�g8��'����O����U麐�r�V^e71����w�jI6��Z������}U9���i�7�t�=���H��`�l�\�}ww�Z�I�'`�x�o'�٨�.q��#�;�q��#ŶO1�h�~yd�*m��Q?�6�5�i��u�:k���q��S�ѿt0'��A��i50_��J4�T�LݹshuWMpn����F�(�?����0����GC=sઃw�a����@�h{���k	/�tE��[V�P��Q����0��\e{����t^�e�Ѧ�p�R�\z\vo��� 1@p�n$���x\����e�˻��l Ā����A�i��D2J��]��#�} ��+ϥ�Vv��h-YSTI�h]���e;;����ߤ���.�9�ת����T��H����@�(�A���,= ������>�`:�5�9'/��J����y�sg�0w�586�g0�@�u3�'�t�����DO���Hk��kw7�� ���?YG���(�ue�P�Î5ߨS/��Q�1��e���]�-���%��`���j��Mc�f�s������.��*Z#��9�����֑ ��xvz]�i���)��[������h�S�+x�w���&}[�T��0�!дylurH)��"6/��A�U0��/�W���[�)�,��H {o�e���q� h'���1$AV����V	O��C�H� ��Σ����]@9V��g}�Y��x{鱭i�(��I�-���X�x��~�5-,��)�V�"���5�a�ZFj^�}�)Q��e@e�*�5׏�q^k"Rp{^[g���x� 3�ο&�������M�o�*��:��p��^�t����\lj�w黍۵����g��z����Gbp����H.Յ�l֥�K�4*g����yuQ%Q;H�y{�FA�K�T)��.�7�k�g�|[<�/+���;\	5�)"i��.Ԣ��L�p23��|�ǃ��콸S�����ގ�Rj�e����\ʦ���>��
S�|�&t-�^��aIbY�+_���	6fh��u�h�ˈi��~�\�E�5�V�.g(��)�������GcaO�^a�g��1�t�����F%��κCP�\O�?{��&o3Z(�w���e*�H��Au"�c�<�T<Z���%w+�3�?���MJ�6%��]���\�x�����i]-9�{�{z/�w-��S��؈p/�dM��/�h����uV���e�����@�[R����.��2m_V�������.=
B�oe�'�p�������(<��u����o��	�Lq�f}s�p�Cr�}`�f_�,V�$\�|��@����f6N�.�s�d�=�u��֠����s�N��ĵ1��Z���p��ý�6�X������TEu8��?�;X� ������U�7^����luU�B<@�lS��l�@p�k�/8�6S>�ٲˬ��u�{�{a�n{_�ڢ>��Z!v>ؓOqݾ^��K;>&�#z�	�J`~Ȣ�pVf�/�}f��f��$
����(�/47N}���,��=�nR[7}� P-�u|v~�����1Si�Y���=R�����͌3�g���5�U���8�����E���g�(��M� 0��+7�i���_^���s���]��᪼-�D!W��3����<*%b�����F#�,�Qp�P�'���eO�8.�����cjs�Km�eώ�/�=���4��ma�qN���Tkv�X�x?^ڟ�fe�(�!����*��FvrgCIġ�%�u����%�((���5V&_m��)�4+�SArx�����L�\��N�ѷ�d斍�b���y��<�[O��a�yU-�+COr��� 6<ݮ<@�tSLY9�+vĞ)]}�+@��"t�ӿ�rԣx*��2�\İ?��_ES�v?�e���Y������L˖.��IYi7N�G�B��\6���po��Wtg=ö��D!偖�T�A��o�t�$v����`� �O3���V�<rn<U���UJ�џ�?�}C�7��D	��ҨU2&�p�*ؕJW��2�*�g�ϕnO��
0��Ǝ�9�#�k�n�0���_m��p�OcG��<��	��3c;�)ߨ?��>j�����C�5�|��[��6|A���N�@.�D|ń��o<��V��X��/~�,%�p����b�j}n����F�N�e����i��B�xsX|ր�f�2�@�މ׼��H���-����Gx�۱�2�h�����t��ݲ,d���������ٍ��[����"����%a��`H8��]��ء#��@��Ȯ5��y�bF~�z|��f�ö�|��g���N��B��'?l[YU,�-k]���޲�{�>"=�i/�X��\y<���1��rt����tEF��tU����j��̫w��KC=�>#|W�Y�� �e�j��\JZ�O[ȕ�'�Tg���{q:M��975���B��8\^��-O{��wp@�|��Y���<��L�c�7��t�g��Զ?e��2���(�:'ѣ�?�Ԛ��ћ�v�y�ԛ�g���c��P������_��9pht@%R��~/��XK������aB=?��`�M̘��p��������1� �1L��$#��B��:T5��~\��G�F*�E���7���s �:/m���{�|dM�P��&��YhЎje�$y�&g��)���@8)�����bmQA�7j}�9�ǤZ,E�(�pkh��VHQ�Pk$���zJǕVn"�Uly�� L��gϴ�o{���43l�r�C*��4��4_���Pq�:%��PJI��7y�.�NucV/j�Q�g<�ft��MML$�i	�N�$���`��d��5��}�.���p�i}�-!Q��t a@sG�nSV��&�E��m���Ty�&�Z��ZWH�_r�����L��q@�U����b�6��6a��\HHT|aƪN�YƇ�8��'Ǆ
������mƲИ�_��2��Ekq\k��:���l������M��� �����Ч��!�Րύ���d����*��6���������o��|�>��S >�^��:�S�*2��{�ds#���"��7CL��ݒR��uS`b�xX�������c�)���e1N�!�9l|��g.SM�2����(��D)��>�O��`3�-Gl�=��K1Z͑?oDf?Q�I)�OL�c1��g��'[�< QAT��l�R�2`B������Y��0�˔#��m�� K�Ailb�{��}R�&!�b��vmPt�c���@	u0K��Ȝ/G٥��xK�:���!\Ut���x��Rn��ze�/8$��e�Oك�LsKl[��H����[2��G�x�Ҏ���aG��B;�&/���D�����W�wB,߮6>�5��r��!��~;�ۘ$]��������I�[J��"݅Gk�;¦\�K$��Sve�M��مuܙ��.p�e�A�a�m����8�QI���z��Zw�cI���M��Y6�;�����f�z�n`���筝�V��������o��.�TD �=�V�t�������;l�.>Ԡ�!��Xu�S���[�V�Yй$.V��G63�~�L�k5��ǭ�ȥ�����2���v	�/<��R&\k���	/_=K�gc~��H��/^(���G�׶�M�+_�ͰU��&��='f���.�HMK8aeC�-��t`9��r�t�c�c��������H�����2BEE��\ΘUq�H#���qEeBMyQ�Q�B^���u2�l�D*%f[���e�W�ė[����ބ��w�^ ������� �Qؽ\�yIOxY��W�@P �H�8�q�;�3��G�7���*=�5	@�l�Pg4����8ރ�d1e�IIM��zs=K�h��!0޻��P��x���4���+D=��=�G0c��4�r֭���3ml/����i���㯹n��n ~�1uݡS-OQe1MS/��Q���s1΀1�5�9���!� C�9V�Jh���G?G'��BR0;{�B�����Yp��n�c�%Bl���$��ᣤ���	< ��ܻ'�[�`�o} L$�hk|rHt�����=I-��\�~E�S��l�ߞ��@){vm�y�F�U�6��@�W��ɇ��պ��"	/ 8895�i&��S`HD��v������@��T�
�Ƴ�{�:��khi�1Ӽ��|����>\T��,�z�䮅)<�Q�@�@W���k���ܭ��z��n^�o��C`{*���xS,��軑��Z�a}�����P`V���µj�Jb�:V���	���;�(z
���`�[0~(�.��`�eQ}W^�X��kp=�'<��>i��_�rL�J���(�0�?���*^����\��b�`�/,�=����os��"<D�ތ癣ݭ����Z��Q��`�2�}mu5�a��P�X�	��RV��
i�ͪ6:|���8��1�Q2V��QW�'Mɼ��r�Z�OZ)=s�W��R��#h@�m:ѫ��j���<�� z�A/[����<����믅--�i�!��hvRRrb���K�M�.�T��� +�7��A���������q`-���)�n��*+�=r�m��꟪U1��i��hw���7�U���a;!1��'DO���E��*o�B�RT��������̏ �(����d�H�K.�ߖ��O.,��8ߎ��U�W2V933�	�	�-6���ϓ�)��(�kߔ/�n�ųHSgI{�ǉ�������˃//p��(^O�`m�t�ɿ�|��ΰ5���傔��3&G�_�E�\�G]<�}�=l3���>h�zF�����_�ȥG=�D=Ѽ�IF:��ຏ�i�UdJ%xz��W�����9�Dv���t��в'ɒ�����7�=��j�|T�op�D/�"���)q��-t�{Upѫ��;#��q�삑���RA�Hhr/|� ���`џ�7`�,�.���WJ���`�υR��;r������Q�����AXm�\�b0�S0������9��a���b^
%��."�:��	��r�C�	rD���ꝸ<����#�Ǯ��fGzerEOF�v(�$Œ��U��f_�q��sB�u�-�.O��/&?8:��E��BMIX��H'�e�|�]����Ħ�/H�S�٧��V�l�/��y5�sq��j�he��݌/��y��Iӕeo� ����1���gk[F���c���q�2��9��K�̅4N�ݭ�ƪ,�M�.�M��b5��/%A�y,��wGV�{,�GКD��-�&-M�.��n<��hv2��\|XX��Z�A����9-bxxx	<E\5� �ڲ�OD�^ť'��Ȧ���"p��x[�[���˲ӭz�C܃:�ٵHх��^�<���0+�56�E/�D��Ũ��8���*`0 ��̃i���ϰ���bb�+&�:�Y�U���LMMkڙ
E_��'�Ƿ�0���Ɣj��W#|����(�
N��A�=-�e�A��>>=�N>0>���H����v�V��	��0Z�$*�|��f�ZYY!N��w�	u�X�."|%�YZG5�F�hG>-T�Q��uwu��V�}�J���;���م߼�h����өY�9�*='?�V��%P(T�ULJ
<P�:11�[�_���?��0^��>�k��6RY��	���y��y��G�x������u$�7��kqU�p�ş0J�2<�^�nh�	;zӐ���=�n����.P��TǷoy���7!����d�k�]g�`��B��d���Z�qh��X^�� ��'�b1Ñ��a|$��lCԝԟ�OM�?;�\1_�b���j^7jd�N�y �-���x�A��M�d�zhϡ�9Ɵ��ADh�k�CZ�hj�v�Z��χ��q�=
,����������L�2˃XyM�8(G �eB�ج�o|��8謼���w�kz�����[7-�3�%�r�s�l�KP��_m6�ub>o7�
��#�Z�7hU��<�'D*R��]ID-����]��B�6%	�iw��}۲��� nn�&����f��D�������e�\j�ty��[�Φ)�ܪ�:�,�}��L�P����zY�c�ɥ.z�P�H�����x�#�������}=-44>��_FDn�6N��ʹ8Vv���� V8,��H��J.� ���|�g�5ӬH���mJ�WX�}��6̸�aFk��}�o��FE���H�B��Qsp�[��h[���e<骎!!�%��v���n�g�qjמ���/|� 'i�#��8��nG�`S[/]�E�$��']^��Lzw˥���z!ºa2W!;����~G��O=�����?}@��	Y�27\<�%¢Rv���e0�9��B�]��\����.ZLwE�c�D'��B�8F�}��{�F��g��Jey��Y����l��}GV��uq�'�G����PݕOW��:����G����R��T��=��kG�$�&&JZ{.v*${�{I��S�ӄ2'/�NWRSJ��;�A�g���ݨ-�����y�y���g���
%��R�@����U��z�f�9�����#j:����e㌲������9>i���7�z�=���_��p毒E������f�T��w���a�G5������CN��D=�����g����f���_��}yX���1!�95�3o���_�b'<MWfh'��-�y/�ԴC����af��s���R���>׫�x;�>(,�u7<P�д�1��[:!!�݉苎��/��۪��4mu��l�I���)�}xϤ�۸�.��d�Yt���td`#W���Q*k��X"�`�J������M�d*#uK>����rb�3&* ���)v(���fW�݆�����=WiIt��w18� �`OS�J(V����$�,11Q� �����&�fACv�|���p����l�~��Q��@C#����s64�Pr�������{l�s˔[ �����ZxΈ��L�ݦ�$��h������|g��ǒ��@:q�����n������}��#����=�UV�� ���Y󈉿J��8���$�����4�H�	�hD��v
�/�^;\ }X��N����\7�z�����<P��`���Y�
���iH�98��[O�ݾo;1��	\)Ml	��sp�[Òz�\�'Xt��#җ%S�b����6f�>��uu�tŦ�ݶ����mW{qo=�༴��2h�׷<��&�S�;:4eh	1�*ߪ﹌��\��lͺ��)z��0�w;�Vm$ ���Q3�p�ƥ��o�1����9�����K�c����Q�v��2%Ie�tl7���\���B7 ��a�?�!�a������ٖ�P��8����|�
���1=ey��#�%��O�p���)^f�+L�
��t��.�� ���
p].�L��f�{0�ż��@[�`���(DN%'>�;ʵ�?��.���LBЄ�����C|�t� ���H8���-l���x�B���s����>�)CS�O��#P�y䢧ݨɻ�'"��3��� $�|MHXrn��ˢw\��!Q�=2E��7%e�z�q�jr~�g��.���a�����Z����>���:D옟@_�n`OJO��z��	eD��A6�9�*C1�o���G��W��3�w������U�G�^���)f⤭�<�\xǦ�[��B��^pD����7�k�!b�/KA�_�^m��1y~x���KF�-�g��ٍ��������Є���I$Ȩ��P+�q��S��D�m���h�Ք�@ ��\��{0�Ii�Y)��sTx<�l�A��DS�g�}�o��~~hHy����/�(N�0��x�0�O{���9���@&s��i�H��I���)b#3�M�/�����w�}�D5�8k��z����u=%�u;��o}��%vrŢk��7/������_�y���Jּ�b���(.4���l�(��U���6�~��4�'�E�|}���d|��X�R7��lD�׊�nO�ybY���vBd'��mB�@ߔ"V�-sel�Zk*S[��h.IG���ąc�KT3ڴ�Q��jWrB4�c5*�N���o��I�D�>��״�?\����V���
�h�M�r�)�8����Ѣ��Ngۘ�$��$�PK�n?���C}��7@�^XL���
�=_�Zp��P�hA#N3��@<���9E{#C��I�"����v8���9�UD��<j�EeX��=����yl��L�~�z�7ڬ@���A����4�i7;�6VO?��7P=�� ��zB���5�m՘g�)M���|�l�շ��L 2������ax�V����>��>}J~�/��J"��#/"_[���@�� ~�rk��K���i���iưe:��?��X�`T)���Hm���s��; �k���!Oc(�����zb���+ybl�?��'4:tc(�s?��ٚ�|��cv���H�~������\�kg��Mڮ3	��>Ҿ�~��kKI�E��.�M��@Ko�e{�Jj2� �վ0�P�?Sd�+[FS�͡ՙu�a�!?���7(Ȓ8������K��x[^��o�o=u]?R�������V����U+�a��3�gJ��D�]5��GS3jF7�`lf���uH�Q���K*x�
C~]O�܅]�z��F�kp�ff�?�b�F��
� 7E|�7��1�@�	�C՚�q2vU�F���<�U�t���a��Ǆ��s����2ɀ����2��7��]�!�+o����S㍉� �''�<��k�_��U�%�`~��cgSŗG�0�/�u�t�3p��49m㊿"T�9����2�q��Κ�}��T���e�C��N�Qr6�nM��<w��eLp��z��
��I���{8��l}z ���3	�n�(�1@���3�u�[s�~I���􌱦�)�L�����@��ܴ�|�Y{��|}}�����5d3K�u�7�����/G1��5��@��_��5���^ღ�W��+C���Su�Zz;9n}y����:�W����8C��;�n�?�u����������d_G���Y��������w�k�w��V���wH�Y�Z�#g��;�*�L ߣ^����l�O�D4ey٩߉D�����В��%[��BsV�뚬 �q'��C�(��_����g�bʟO�q(�^okl��C>��4ט��x1l��^7u�vwݤ�C�;�Y����I���p/��4�@T1·]]��}6P��[�1�z�ű6}gT��Br���j=}�B���M�Ok>�_<���O���%%%)��LE��7�G����ݺ�ļV"�y�O����6wv���-�m��hXk-M�B�������ML��Jl��$v��<;F���Ӈ�,��bs��}�D6?*я�jI��Ե�RYI�/��� ���u���d��xe�X��e�;Q0������-�^	E���;���:���5��ıWYf�J]�M9V�\L�L%�������?Z^�O�_�q��ʗ
n�\V�������s��]W��.�ض�i���8�N�9m�>�������I ��Q(�x�y�s��t>���t����K��� S+x8x���u���o������X;E��1����h�Y�$�ϭ];��>�	@�C����EӺ�֙wh���.�]���T��B�V�H�i�����H��wO�ۗ� x� ���n���w�&�<y!��c��)Z��x�q �S�x�2��_u�-��iwX���27H��$ ���\q%�U�xۑV���8�t�%�10�E*Đ1����J�6G㵤gn���6��B����� >�=;�
�N�)�Fه[p��!�V��V�tL�{�kGW�/f��{rc+°�C'++Y�`� �8�����?�Fp�)�d��#,f����������8IKK�ى�

�f��9�+�G6���4`����Ht`
��d�Ϛ����E	JJ֚�����Tz�6�Ԓ:L�����{ ts����=[t��{�U11�D;��J-�C��t�!'�}n=G��)ˋt�㶑�8�:�S���^w�\;\{���V(z5�
=�@�\�#e� 47�C�Rb$� rc�7g����F�ͦt8fN��u_>�"��yQp�x��Ծ�mӖY"Yg$���n�\�<�'*Z������P"�`N�,��F穲��5��#ז�����D�kh��WoW��몖����o3pi���M�?^�W�08O C�ı�ݵ�q��췇�M^�;f���{���d���a]nݧv�^b��o��UF��BEGI)���b���4� ϰkS��ݲ߃G%*U�G�
��Tj5�t��zJ�ޔ���z�$~zL� v� 55j@�4�t75�^?�9ܲ�j�.��ދ���0e8�K8�p���%�;~N�p��Uw5���r��p�ȿ�|{��\JUT��5�K�Ąu��wBC�^g����fU���.R�i�_�N�^4��O������͗��k�l�Sq�V����i[�_�7z������z���w*���+MdG�gO_u�b%�<�꺱N��F�螣G�@P i+��@I�1%y�=H�������Z�7�2L�.��2��g���n�T=,t�-!f?)3�uY�t�R�9���ԝ۞��8 �a%@B]Nc����h
�g`���J;�Qnnl���/T�&��4�e|�;�+��2A�w|�q���i�Y-+-� hkر[z�:��I�9LU맔κuh�\�Y
��t�����V�E���>Mڟ�y*�^�/�h��׼�p�}�ۀ����ŵ������ͻ]��������R�?)(�����+2I���O- z�(���iMXZz}]�����~š���&4�H\0��CUM[�C[�����=�`�/i������������2�_��Z���7�7qڧBi�ox�O/1����>�uW����wo�il�}J�X�{y5X��M1��������~[��d��MIOQ�ǥ%�L�Ώ�ф|? \�"��qV`c��OVC	�sQ�ǗkQ�;q �Ŏ1_�[�:�GNn��ϟ�3����$ Q�s�?`E%�)൮#��MRw>K�Ի�K����5U�!�OK�J#�Ȫ+�a��Q��#� �w��m��+���/oX*��2
��O�.}
qt��L���\�E���X`�o�i��������QQ�_��H���� �݈ H7H�tw�4�-=H��R�]24Hw�=�����X��5Xp���|���{i�;���c�.��n���,Ro�J�fk-��J�m_G�8P:�+�k��0
��z�D���cn	�z[q`ٽ��tH�����ڔ��/t�{0�,�=�Ck ��n�H>������:��ѻ��w��7ʪ��'����h���e7�tyqO�C׼p]�v2��R�y����������511����$�ˈ�i���ƻw���,�|��,<=S�I�|�������N���3Hm��6���}i� ������G�W=$\2$x�#��J`{��N:ۃgX�>��HY�׀ԟh��WYë�hP���j�!��<�m}ML�e��gy���*�z�]�;O�M�!Ȫ���Ի�yf�l�	���,��9]s��ۓ�X�-�Ow�jV����}�y�U��D0Qe���8n܊L�\~C���?� v������6"�	pa���������?�3���X8�O$R!E���V%M��;3�7�_�k%�p�.�﫯�K�'ةUe���~��q���b�z7X�J�VU9~>��x<�\��\�L�ч
��h�ri@����a������pY������ZU�0��sK�A�=�����Ő�H T��! ����� *�-����OOmmЯ�ƺ�Sv����V��|�����uR�k���m�4�b�!9EDY���J�(�z���S3@1�lK��E9.�����];[69�����p��Bm�����r���Ђ~f��;%\��Es�OF�A�����b�,SL�i=�i���eqs_���(��g���(���Fb��3�=X��O�LYC!���lOP��Z��83��l�2�8Q:i4���2����<a��VO���.����&+���"s�N\
UG�S��݋wR�m����㬭jj�y����+���\�*�Se]��A/H�r������ĺG�B	d�A8��c21YGxn����P��Sl#�px��5�/8�ٔk;TH����������]��:��Ǜ¤�16ğ��4��W���E��vaT���B���j��H�>����=|��jjv���#I��Q+�n\�j�TWm�4J�+���?U1lL�d��.? ��j���	��o1%0^e�u�����o�>��b�H.�ߓ��=�6N�� � �Ι�ݯY��Ϯ��q�ekN3*��a1_��KMÃ��LS���*��dBv��p�n'������5��`�2_����B�[��y�ns���v���ߢV���e�D���~�����&����d����>y���q�� 1�g��ƸV��tQV���:����n�Z$s�s�k.gb�^�[�h�5���f�n��o�W�)�:D�T�o��l{��n\�z�&�眪��Sĺϱ��3���s3w��㚿�%4g��]�=X����|�t�j��5��`�PQ�͉�Ԃ��Z�¡�b'+NΟ[��uC��'r�c*l�		��M����
)�����J����US�	�dZs�c��^<��c~gyh:K�J52��dԐ�д�����V�pv	$bpP��� ��pƗ2l\Q�����+�L3 ~RǏ��h��t4��Ŧ]O�lQAC�,�16U����K"�?�ų�yb�۾�n����YD�6Ɖ���;���A<�_4�J�2����O�]���-X���c��R�Z��/R�Az��lߌ3��������4B<��3�;}��4R���T�ux��5�"�'*#^O�g�7B��׆�/z�>�������@4�p�@~�8l�L�)2�q�DE�Ţ��'ϡW��U�|F�UQ�oP���ob�S���c]���ը��m�X\��Ax���'�?*��f{>�\��;�t��Yƾ�����$����!��]1P��3l�Bz�&$$?�ۙ�}U�$Ϝ�r�r_Ub�C6�'"eS��T�T�id+���w//���_zm������/��Z���v�j/��Ч�C�(5�5��yƦ��UoN�5Ky�]5n.N�mOw	�������6Aq���s����
�mE��5��G�>e\���Y	Fe	�w�%��`�����7��iD�|�\���>����*�A
��-���G��O��B ��@W���9�o�'t<;�E�:I���q^�4�.����w�1bQ��9
� SX��{�/�F�s�"�&��������qr]�+Wttt;oN�N�ZX�8e��C�ɨ+F�w�f�0�qk�Ӳ�1f��^��e�% ���WK����o����F���	� �9QҩS��9�;o!ӿh'\<�$j���ג�:;��5�>��_��s?���̆#���ߠ����G����"Shf0�ve�^���S�Y+�*4s=�0{B��dD��_�(�T4�PĐ�YurJJ�����BLL�
n���
&h��.F���rIF�jt��=�C�ʾ4��:����Ҥ���C��ސ��;'�c�p��]��R"RR߾�!�j��	���Y푩u�X�G{����{�,J���hk���.���������8��֖o��\��
��+������QZrϣm�^<?l'�0��Q���n%s��!"W�"��M����Gc��Y���{WBֽ�&
0�J��ތH�2\��`�X��n�[ėR"��|Q �P�H(��7ˢ2D^T�\W3��/�}����-)r5��2>~	s[�Xӿ31����p����z��>(����6����v-5�tA�V��G��("a�G���t�G�K	g��%$��E��=K@��{���TTt�+��!�VFg��1>;�.N
E�T
�K7�=��q&b
�l�u�"��}��>#{�<Z57!����н���t�Jw��ۖ������U�'n�il�ET�� �������Ky��~^�����ϒd>x"w�1�n�z;s�� V��"��"�5�J��i(�q�ˁE���/�Q���K�_��K*(`�2�44�#{��w�����u��S��_�vz��ccc2w��b��a���"��I����/&=��'�5�]���:���
VJ�o�"�Wn.�/:Dn:L��+?kNp9"gH	;�!��)+�)�2��w}�I~fS�թ�A�����s~�ޙ���J��#����FB�OE�����9�_8K�^�9�޳���\z��sً�&X��ћ`	@"��������Y��#��
���[9q��&�u�Rd�_'M��c�;��4ajj
{|��ѡ�h�Kc�ڀ<Gv�.�Z�>v!��B���|xl�ӑ�l�".���	�t�%S�;eJ���ĜI���NQ��K�+�ٮ�z'ۤ���o��)�}�/:c�U��ĄC����uCƻXt��"�y=�w_ J����v}���~����Z/�AdNgˑ�[K[,'ҏ�w��~���\�� ��C�6�7����^���M��ԡ���iHL�b,�\I����K̟�q�"ݮ�7��=�b�v�D�0 �GҎ.��V\_�{�͘U���R� >?���$Q<�<�G�7��8l����ˋ��\�>��Ҏ�+��y��)<�H
�:\}��F*ɹ���uJ3F��9v���F�֪~~��s��g����C�:\���>JK)4����q0<:�n�eʀ���L�#��j�A��E�B��L�mR1�a�S�wT��{����ɚ��Z}�z�@��c�X�pJ�V��ML���r�VDU�.)i�h������^�������׭O����B���\��1"��R$N�J_���ȊEGw�_M	�u�ϛGh��.��E�b"ަ�;�y*���"]��!��ၛ����ʈ�O������;���6i����OTp���@��5��y���N��?ے��k�	�)N;;y��D�,�5z;��^U��N��_�M�Et����q��i��|��e?5LEN�c.��_fF�5
i�0e,��)��BTD$C]�a�l:x�ͧ
3�X.k�#��	,���D�c�첅'������"�Ps��{�}�ފ�nӋ	#A�5�Q�m⓬�3�D�i��J� �!�G�w����6��x����|��^9�h�~.�=�������KӏÛ���2����Dz��w�r����Gk�G� �����0&���+�0��.�l���I��s�FNV1����`U��h�����p��M�B����@���V΋���f|f�o���?Ǆ.γ�n��2�y��OuU�ڳ}&ː3d�E`	}^��ó�}r�>N'�7؍���x��]�l�}@��7��I�lez��i�f:\ѯNk|8�O&%]�PL%�$��Nj���®F��
�w��.�~ɉ6+�����\1f�c��]��\+�˰`����l�̢7c(A�4^��n�i�~=�01I:5Xe�$�ڦR��~�C��݊%n�d$�ٸ$c����U�.����o���Om�0y��~�Y[�ȋp�4B��a?��Y�?�z��~�n��?�}���弯/�60F�sI�O���E���/~��o�{	��`ϻ���^�ę5�@����	Cb���CE�]?>E=d��c\P�hr^��������/�b6,W+0_
_��{��'�<�e����U�?�mʦc�/��9�p���uzk�˥�2�«�����*���"�qY���Ƚ(�+g{��6�ܿW�9>"�5��+d���~zU�'�#4TȆ�\$|<��G�M��|g�P�����2��czD~���1�W�(���]�����3�J`m���2D�����S�scp�D��2�& ڡ���k��������
�E.zx����s�5s�f����v-'���W�c�g�-���v��a�A
ގ�w���kA�
5��Dl��7W��w筧'��7w��V��=>����{��#n0-z���[|x��𘅸��\���c��ӋlE��-|9,!��G�
�X��+Gهm��\)9�>��@��z��Z�6��H}U�o��_DtR2�9�^*Ȯ�g�Ǽ�@a�\��z���#�c:����A��N��� W��h�)�����r�h�RS+_��U�Uj��:2j�d�/��4��a3����:l>q����
xB�G׏/�c �_�ίs,&�VX1���f�	Rd����5���;ׄ�q*/G����Z���h�B�l6, ��'�5�H|D�U���R{����5Ƞ�����u6�qC�Ƽ�窢���������+�q4g����(�Vjb���5��ev����?4�:A:G���悼	�����w.���棍T�~���q��1~\"2R �/�~�5�Ԝ0lz�y��G� m��K�i� w�K��^.�AJx��#Q��]��'��%�+צ1?CbE4wx}+�&>��HQ�-��o�89#�sgǺ3WD�#B���U/�SY*B��-�*���!B�}�:ZC��%*�W)*��z����䴴^m9c鋝���:����A|�n\8]�7��qZٳ��_؋̏h�T�%& �E�rp7�(�"X�1>�*�Z$��R���#YɨB�ƥ�)��c+�tZ����_5^;����f6k�����܌��H��>�^�::k������'ZkST̖�	t���<�hqb8@WW5�d!K���lH� �7-��r���'T��z�����r+9M0~)�
:h�>[�G������{�J���TIWW������2\$-����B˯�ηߞ�/�6�%��󅉡�ll.��p��׏s�˱���.'���m����#��'��A�HY,���.�]�P��Ȟ�0)nlF��ٓZ|7�l���#h�t��uk^��aP���)\z��XO��,����yv��׫~�Z�h�H�����v]�F\>�嶛�b>^�zj�����A_"3��"��`|lj�'��@\�x'mK
��a�o����Tgg2+�@6������1��łW��5w�XЋ�X�Mܤ.xT`��l:r�utE���v[+���[�{c�uo���������KՌ�׏U�ʦ(RR-���X���d��_C�'ss����>�,׷D��bff4�_��"���l�oT��eoi5�����&�]�����6F�&��C8��(�D�S~r$	���������]�A/��X����G�zu����D�2R��J�c��kw5iԀ��h�j5��W�o0}�ND�ד���U�������W�̇i2Bw"w]�PH��B`c�MU7Y��4� E2TI##���+�7VO���X�:u�)h=����鮪������2�/5}c��*;�X5��ev��as��/-P�ְ��5�����;侓i[$c\�urv�\�פ����2޻��As��{���9	� 0r;���:���D����iY?~�w Ʀ�N�¢�u�<�j�H�'�lCՖ�����g��|��ࠧ�?4	%VVV{9�����L&%r�e�8��H#�v��R�-�S���g��d38��ߖ��8qCmS
�ݥܔi�1{xYY�g�dM�����s�J������(�Q�����z=V
�"�ok}�[!��_C������t|y���3��N�b��"�adg*��.֦���궻�'D鑹�=e��D8�^��状������_S�;��e	�wգ�H�}Yi��@�6�<�������*�./��6 ^־�Pe�Ƙ����At�S?� ��7���*�!�y5=[�F�\T_?l�a�QJ��
#6�����pu]t�/��)��(�1hZ*�sg�˩@SM���S�yjH@ \: V�INcg��_ޯ}�%~.'��x���v1�_�f���.|�פ]�lw�.��>�����?�H�W=�����X���~%�Y��W�gb6e+'J��P]天{)۾������#\3]h?b���K/�X�5�l������Lu#:�H�:��W��ل��m�����Ϣ��k���﷪Dx8g7�O��x�
7'�3�:W��`JD�dݕ�(0f�F�f�����hc7��G"9ش�JW���?��#���?3Q��ظt|	��{���a��#��H� QfF:�w6���o��6Z�rE�*P|�o� 3iLn>ЖF1���%1@tF_�RƓ��?й������'9qY�@�(<��:�����=��9�غQν�ڛ��5Zy� ^�`���_�b��v-�������W�j�ou�2�q��hf�s(����p��ʫ����}��h֧�f�zkgǂ'���I,�vv��w���x۝��Ү_ ���Ct���`�/>|�^��	�Wo߾@e)S$|�U��|��Ƴ�gE �[��5�/7f�;5����&!!�k7v��d���":#@�2B@�P��i��!�]WJoػ���9�%'Һ}��42��k�4;Q�6AJ�H��򾖩]6�RT/�]Hj�BAIU	�r�A�@�N��(Sd������P�]]�k2~�3���_��L-x����`5��q~���h���F����b��<���gg��aj}��"�B�M�ڂכm�2	Ȍ� �"O�m�M0�	�R>G5�.��z�w�L0<)=�䯨!�}����Ԍ��Ы��E������81�8��p�t� ���Zy�x0��w�8�Ԙ�qqh�g��M��]�K?�ڔ��V���5����|����{MM�Yfy�sx R}pN��Ki�|�ϖy�[�qjjj�?F� ��I�õ��6�G��]}{�)�?�����ʿ�"D�Z^����[�e`��l(#:j��1�ȼ��ڭ�+M#�/�ܹ���坑<����%�u���s��MHϐk���^ �K����禷4"kR"ᚅ~PG5�|q�ٵ:��h؁Kn�x`��׍&Y�9�L�'g_CH�:5L�4��2�e�xz�\�1��TX_�	wN�Ӎ���ߌ�E�t$�;��@ԡ�r-/��^�ϸ���z�8Y����T��5����{��e��ܭ ��F;;�-dK�V�̚�(��-�A�Vu?�
[a5c��fh�0��Fq��(���0�y/�_b�8%���~c)��E�]_q���g�}i/�l�y�$��� �ky�7�5�:j��k�!��"�H�הo]7˃)Ajc�'2%�Ǔ�3������+�1DE�|6���㚅&4Y;2�'�!�$�Z��0~r]�]�kDRΤ
��v�t��G�z"��<;9Ǧ��=2@���Ҵ���jE�KPH��6�K�uTw��D��%F[gR���%5���fa��~`G�=��r�����="Y<dھ��kV��Q�{�4}�r��"ML�����ҏ��pF_=�.0#��5Z]|E�� %?�c�1�����=�6T���]E]1��M�`h�)��t����;l��ݳ�4k�����0;&�w���Q�d����7-�[zܜs�3�1��MO$��<L�r1c��T�\u}�@����,��U{bgܹz(�\a����a"Z�s]����dh�b��[q`���X��W8�u���Ӈ~��Xx��Ժ��A�%t	��(�9�\��8��ޔ`�Z�D�a X���w+��""��G O/�JTJz�J��p_7HЋyבb���(���c���۽�cX?�Ci�ٳ��A�}7�oL���C�}﮲���',B���-�,���������'
.��a�J�[�-4�d����aA$54Ԩ�\�B�8He��tb����kr��U�;x�K�y4�}��e�Z�xy9l��!?$�t�$�$=Z��d��_۱j�c.n��0l�{B�����PR����B8����-w��C�c�w�?|�6It�\�n���#���:���|��(�3�b�Ю��wY[rսYUWR[��A�vu'�_M5-�|�;�gh�?�����yuf7Đ<!��0_�Ȟ[t�g�w�q�vrZ��#��!Q��m�YO~����ֱU��5{&��!������+�(#xA�Mw���8Q��`#�{8۔7�:�HR������Uｆ~�!�߸��w�e~����	�T{8ʗ�/�ł�x3�Vt�Nmi���ô���$$�(��/ϰ~Rǅ���/l%�F�|�T��tk��\�D_𘛳���c1��Z^hh��e�;/��H��j�����܏�֕�s��wW���w�[o2�K�ھ��tҎ�L�9�ϖi秋��{�����K-n��y�L���d�8��[���v������9��þ��!�c��*zI�Ym�nw�J�tuZ�?Er��~g�2�L���>�`��{����1[��0d�n�ϗ�W_y�Z��SE!�o���v�yTz$�?M�N�hV�$���U����8�-�������y�}�Dj�Rh�.����%���N}3�c~'�wr�8��2mY����������濲��O�J����^�6�*�>품�=��(����z���L� I��	���`dܣ��f��w�*���,�.o!6�(� w���;�f�r>>~�w����Ǜ�u:�P������pwe/�����_�䛱,�,��5��j��ɺ��x�pa_����T�$�1w���]���e�tr��U(��3vJ�&-Gę��� W��}�sњEV�5�p�i^��5��hnqm��l�K���ϧa3��{�lpim��l��LA	�H���v��jԿ^�DL�Ǝ�̰�b,е$��j8-��T݂�g����@J�%]����qMJ��;�/�{�2���H@�������C\�m�{�?\�G��P�B�}�_e��w8.�e�7~��`b@�4���o���P�}�i���XѬ�^w�}�j��L+��o^�\�
�G�s���(��H��퀐l>(L���Uw24������b��tĽ��K�_taPy���جLe	���b_s��?�a�߱'޿?��K�oЍx=��Kv�Ɓ��4��P�L﾿"�a�$�1X��^��M��Q^u�bVFS��t��n��1�[�vU��Κ�{,��=��yq������Ⴂ�|��	�5k�I���&3�4��~>��|]B`�l���8zS��j�����R,�Q �5�̧�B`����am2$q7��:cA�|�:&�g�9���F��6�KIoy���il�EI3�$�G�N�_�y_�������l�d��!�8��*C&���Ve͑v��U`15���Vc=��o'kQ]�zL�֢����<�	3p.�&t����Q�9�S����@r��P��{���w.JΡev� ������d͜��M��|O�v��x�&�h��ͮ.���	��֬Wɿ4�~8#��Hڌhu�}Y[�BҼ� rV�����u�K�.Q�7����Y��`\��I*��b?(?wJ�~J;�~�Xٸ���j�����O�3ow/o]I�7�Ԃ���Q�&S�O'`�
.Z����]�.鋴\���ؗ���`���n-��7un�H�XP?D��-P����v�ц0�)C|]Wdaq�o��p�S���j�;�� �}O������ɸ� {�njY��o�;Q��'�F)�_�Q����B�3�NK�6��G�wϦ����L���������q�E����l�i3�j�ژC�����c����l�瑟�C#迃@�����׳���-�m	%�0��1�~5Ta�Zñ��-�<��;��L�V1y�i U���e�g�"e`�8�o0g��Kbq+jl.��Y����7���pE��;���1��*�.��I�A��%�IZE�ngc�s����Ǥ?�D�ۜ�f7���5�4��S׬-!���t|���̀ϩ�yĹ��5[?���8G���Iş��]xyh�zY�cu}D�Jz��>b�Рv�'\UB#�q��8�`���Z��9ҟ<�׈��u�����-7r+�j����yoq^��l���Y��ۙ����E��SpH�%��+|ks6��� �8��X�4���W��s>��*�����.��n�O��8�ķf���H�[!�϶��NT�d���$�_��ƈ�T�}<쥅h���3�?�5�F��S���fw�� Kg١.s>�g'�si޳�La��7}Θ��� ��y����|�_LOG�x�{�9<JMVa�{$��jⷧd�igxyM�FŎwc�
i�߮�@�ީp��u��Ǆ��Fn
('_�a�9F�������P{��@���'l�YU}L�.��a�]�M�-��K��.�����I�-j���0Q@Gv��ז\r��䞞��p�h[�_�J{;��e����=%����l��Y^9�+	������O<p�s���h6�"�{u�����1�'�ô�G����}]����A�����?>5b���n�[t�~ϊ�������
���dcu����I�e�Ϩ�,n{��U=�'�I���F�E�ȿV��%v^�� �X��օ.�~8CH���|�������ˀ� d^V}� ���כ[#փ]
,)��:ߣ��6�aH��r�_&�����a�2���4�Kc���Hz9eJ>�}4�c�"���0Y*�7���{�n�MXq�9=�-@�VZQR���h�/�{�8D��0�,�uw�P�����Ѥ�)q):�|���ð���	Gyj蓇h��4y2��b𵮐h���I�B�������"�x/ݓa�������Z�k@��Z�G��	�3��k]��0�?�6no��3��l�2�hL=Tk�A]xMf��O�|>��u�Z�%�==\����L �۳H��y�e\u����V+��ǝWBf���^Iu�_�ʃS���J�qQ&�*.�E䁶W�tp
�I_�4yx긃��C������,ѩ�N����5M��9Q������������-��
�@���l���Fr�C_���>5jRR�����XU����阬k�{�ǶR�˓�ۗ��9}�R\���#��,_wʙR�`���;Ƿ�����0u�	�Kcxbx��¹��1����Z���wv���@�[����ġ����O>�T��\�K�=��av���S.�n��%e��P��W���,��S�s�f�B�Tm���N�޾j
Yh�!jk����y$;�o@;;��N{!���
\�u��Uڢ�9o1�T/������ZZ����V�ˁYtX����h&l���@<I7\)$�xʢ�^�vW���=�3����O�a`�w���H(6�����FK8 �C��������'��=���\�OhJ�4�FEq)ԝ/��޾柭\@�gSu�̘��'n,���٤h��W���,6����;�/dFA ���#�\k�혣D��.��U��Cc�5�ARW��Y�=��O�������/������-o���A���H��QNt��^��
��<V�*��a$ �K��ۺ=�X縷��>���v�����o���$	4�pQ�sc�[��qw���ߌ��-�Kj�.���˧�̩Ӛ��B~�2/P��ʗg��!����!}�Ãl�w�j���'�K�=)囜C<���WFng�`.��˃����%��u�ձ?�_�����F���ξX���̝��G������k�K\�lK<Ǫ��r"�A���;��=�S=�.�M���c+0�n���Ka�AvS�G��m�TI����.@�C���䖦�f��k;O���k0'/*��'�K�0������;?�y�qlk�)���k�Mߧ�"��F�9��<jD34n��H�ˀ�*��Q"Z��t+�W�%��63���pѹ����H�K�VM�<C�t�o��Z�墺�
ɧ,�IZ�yET͚P�z ���O�E1/����7$�GVvT�n��F�&�L����@��j����ۢw�&)��pA������SQ1Q���j'EF�g�����o-�����EQ,V��"��vm'ME�F'���{=��w�o�~SZ���x>�+sn���3ܻPB�o,զ�/j�m�d!�t�m�j ����B"�R�<�.y�����>��V���~���̛��8ʬ�U/�AI��?i��x��o��5w�U� C��⻝C���o�qpWRNc:���v�ը>�`�XD�jh��W�V_��NH��b�1�Љd���&�&7D��+�Hݣ�� :Nc�����3&>�e [L��'���@	����K�R2�)�\���g^>U��U���Yr�|���|��ٚ1G�]C�n�D�'��F�@�� �i!�wX���i���)����r 9�F+�#T�h6X�P=��1;��uq>�9#�j�!��kud����;L8�s�&�! ����%�"�Y�B�2	��;��_�fVlu�tŷ�Ǫod�VTl6)��i,�l
Ig�6����k��@���;O�� i��V��-Z����Ih��vd� ��E ��X���-�<C���� !��n���2�߁vf��G���c[�$�3��n����Y�#�����E\{����A�ƴ�������)6��Y�%F���!P�5�K/�p9���l��IG����dc� >�����-��^��~{������r�}�N%��٣���k������w]��('f!%�;z�fCi��N�b�i�_��
�7�k��|/��W�Qn�6�W��;���&8�\�3,�%m��{�˼+D�奷���\����C74m��;���r�[,c-~���.�֓j���F ��t3��gng��-�cZ�uק@��cHjܢ���'}]����I��lV�����e�zNp*i��6�,�S�+*ixMn�!m���I��.��(���^��+��:�ax�[��wx~�_UOz��'�L��/���{@9l��X�<F�����h���/糛��;U<_ۉ���r��� ���5�V���K���3�H��ⲱ0�լ�P��m���{��!������Qjq�$�`�pM�J��/)V�p��2�wH'�����Zal�eA��)=�R1�}K%`�C����6�?�S����ߠ�~�Gb�J��t�c!����$V���n��L<�yxl��)�\���i�U��E[��ʚЪ�d���i���ހ5���N�K�c-�?:� ��KRW�pPU�)v~O@��������M�R<�Lk��t݉�F��nBLA�l��볽��]ܔ-�Np�Y������]Q�Rwᔟ���4M�3е��4a�B��u��Bny�-����/�\�byT�*����	�	�]�tC\Ѩ��a&��;�͸x	��%���w5�������5��W�8p.v���U��[/]旷�N�)������R�u�����t�ұ,o���KX�ͨ�S(�\"��c�n�㯩���ԡXr�tS����eޗ�Β�J��C`_-���%�}f�iRM烤��.{(�J5��	�d#�
�@�ݤʭ��N��Z�A�X	"��cMb�H��dcĽIdt���c���x��Й�|�L�n� �2���WJ�6�~m�#m��p;{c�ǧ��]�{I��y,)�=<� ��-22�i�(��ä=��ܰY����om��@q��ޞ�T]t+#K��v�[��]~�Ud���`�k.�����T�x]��hS��:{9�nA�K+�R>	�eEl�Nu��V�<R�0|"K��q��U?�\�Q5���zb��,��0a�ݭ��5z�#
!I6�����;��{L�k�a�Q25{��e�wH,R�H�D�h�[|	���=%L��jm�����A�'��ҕN}��"�V��a�>2 ��Ҫ��CB��z=�� j���ya�&kR�/ooKm�t0� @�7zDl��l��B�wHF�\L��O��l�Ko1�P�~}HN��}�"�.(Y��W�x5D`���EU��%o�F��f޴  ���y9�#7˫��d�:��g��t��(iZ�`fH^�X�������]K7=Y\��IE]�[��@�Q�@��ŝ&RYJ�6�\�I��X�/jjN�$W��ݺ�/¯17���d;x��D��@���9�t�����A����moF�7�7��b+I�߾^�Z��	hw�=�M�o�B���`�?��茶���h�rH�\p�[�o����ܼU���|�xQIͶ��_EM4t3�7��C3Dr�v�s�����<��n���I��� E�sU�\���3�@x�#�[�b=�-@�2W��-M@@����������})��^����d�ffeZ<��5[g��A�/חlO��<��_<�g�t�̹8�������䊨��\���H#{0)O��
��\lݖn���s�!�\�A���7��)�vj�C��^��\��Ms�f�lr����,��:�H�7a�o{��F �Q#ܟe�aͯ�"��]�?�|�z�>H��=�F�«��O���jR)��GH�����{D�/��Y��J�(���B	��"����^�&|u�Ҫ�	�] ��bi�q;*��|Q���|$�PD[G�E�Ւ��*�z�����͸06�E���q����l�uƎb-Vj��i̬��XX��V<17[�L��mh���9N���uj��5g�Q�J���q���@z�k�
65n4K6M�eҍ%���	G��E�򾫠:`����R9$�'�~u���_�>�>u��ܲ!9�ȩ6ьr�>�&��ۗw������[��\J�ŋ;�w4X�{��}��Y�U6'�L��CP5�#�=�3��$�0�>�O��/�ْN/�=�/I6�9��*��թ0"�kjsY��+��KY�C�AB�❴�73��wܳ���3b~�Q-H��
s<��C�����`�j�u��ؠ��V�^���
�$3�>0�l�/���y���&;��J�֨$CS˪;�� ��]~�d�2��	F0-�Ju����qjrF*�N���qu�]˔Y��)����b��
.��i�r�0���������&��9i_	�Ƀ�J$;9�w ���:�8�Ϝ�үo�u%
4���� @�.�_��+���-[ �6�P�9�,w�I$�C�ԉ�n�)`�"P��r?U�����%����Z��\�ڑ��Q7����<���q��n�hn�}��sF	��mئ��r��] r�xm����NF/�Z���,�ԗV�z�.�K��D_�^����}�T�=�4��er� ������ B�83��B���L�"�0����v�jW1c:�����II�������x�M���FQ��W�����ȱaK��'OE�l8햿N��v�&ŋ���{X�g �����^֨F��F>;����?���}�hK�����آ�yh,��#P�O�����"x��_�[-����(Z���F�t�x�c���He
E�͕�b8��u�ɭ�����*�YW�o�S�y.����N�ʸ9&�ˑP,�H�N�y�>Q��+�����}c��W D�|z��h��!jӨ�����	�-f]�B�X����V�l��]q3���U���^�޺�ٚ�km�f��l��Q'K����=�����Ugꍽqo���$I�e�W�\U�ݐmc�����7�<� ג�2�!x-���_6ate�$uHj�]?ۧ�í�A�A�Z�*��T ���:2@��N�B���,a*
�����a�U��]w�ԯ�iS[�p	���N�:��x)�Ukw��U!`�
��椭�7I87������<��p&!(ե�G���|#M�Э\A����G������z��/i�	��|& �
��/����p"к��^�'į�,Z^�kv�Q��y^uT�����WV�S;���3|w���
֨T��o�Qq�0���`8�_�0hW�����;w�u8f��R��־�����\�ͻ�B�r�e�1�qjer��� q�<�?���x��/>R�[xK��BZ��u,QYb�,Y+��o�0�T^	!d;ٓe��P^�}�i��$�c�0��jy��<���s�s���=�޹���d2uD�y��P�[fVU �/a�rh5#�L4�zE��#0�V�p��L�az���К��!_h���U"������3|��#���
��<��s�_��:��2�n��rʳK��3�Z�C�Ip���Ӓ!rZ�ּ�st��UՄ�w�ӝH�P�;&7���[����%�U�s�~<p�Y�aq
O
]���-��	�<�_�[��m��ßj�V
Q?��q��3>���,9�iL�I��~˸��b����^�Ѵ�����n��/wiZ�{�+<��Xf���j]:�x)�����p��|�Q�q��(��a���:r��i���#vh-0���Ǡ<�:V,�ʀ�#0_7&�����*�q�]�F��r�h�&�����T�����]�u�1�<���2��7�>�{�Ԣ�c&���	w��4�J����G
u&.��M��G����ڎ�6�صZ�EN5�Ϭ�%����)���տ׻��䶴$~�l�޾��m�ꋰ�-�Q*g�<�LX��>�<��m�y��޸���e��]k~~��28��@�m�X%gZ��lp2�x�^s�G��(�ҹ��@�`^
?�?l'�#t7�o��;
~s,c��F�ZWՎ�����3��fX�D�0���������2�fB"���|�5�M���F�����;�0���5u����jaч�����@�4�[r}��a��q��Uy.�R�vˤ�F��N�Bo1wϡ��3}ˌ��}}�ã�;����hR�HE�%��ʔEig&���0�[QͿ�;�W���؉WW�S篇���[yQ�a���}�t[�sY4n�NUU�������L�_/�o�Z�m�.�p�����Ғ�ө�1�,��"���%=w�������t�e�m��V�_�܁gV�)Y�nח���������q$<g'!Ɖ��l(�>U��i��Dm�ٲg*5i6��XLM���E~"�_�E�e��TMl���s5��I<�B�w+��c���<u����V�3�:���Ū������
o{ԕR,��q��-���3��}��8�ޮ�yʪ}��nHt�\�.������#�^�W%��-�n=9 8,&�M����YP���q{`>.�g�8�S��w�ߙ�q��2��򓿰Ar�:���fN�"a�L�Ӄ=#ˋ��D	�c
� "��A?-w���}!#�&#�m)�r�j�[\�)Ύ`�!�2���h;��;M"��-�K��}Y( �H�&���7Bύ��S�V�<'*Y�M�sJ0��F��~G/����^|ǧ���3�FE��ִG��V;k�3�i������C��+#�O�g��y�-��$��
�R������4��v�Nj�{@_ψ�uR��Q)J���>߇���r���K��k��b"Y��Wޟ]�, �j�^�F
�姖�z����殸ڄ���M.��j�`{LC�@L�N�D9>��M�j�M{pK6a'��m7�9�!���E�g5�*��.ÿ́dW����Ry�P��S����_����K�'0������}���<R�"�R�ղ�\�~(�@�c�ϐ�[�Z�Y0��X��`&nmWt�7�)Dy��Qz�0R�q=����:���EL�Q�С�Ɏ
�ӕ�j�*��{��y�ܼ\�e)ߴ���W�U���j5���3������`��\]'G_�G(S��BN�����_�PQl�,;��)���Nr��n�6����:mf�}�Q"+`ݪ����M)���(�nӃ��A9D�Y�%[Mx���鉿 �o4�z��x�1}ϕ���d�:K������v}󋚛�%�%��i�b��;��rЉ=xp���½S �����$�W�0��K�)�(��q�������{�47�V��_��UYc�^��Q��}���G\���e1�c��0�&fͤ�X�s��ۀ�j3��-7�"�(:U���S��U�8~�O}�_������2�mKd�<�D��T�mu�*������ot� _كoA��'��A�ӢsE��!�S���u��[}�X��¥Ԛcjuew0��3�ja���E/����C��c����s�~���{�;�%���k�!�^��<���!Sno��)x�e�,B[���ja���۲Նɪk*n���T�X����1lenͻ%�`&��.�
�VͩpEXv�͘5��/7�}�l�%�;{�q���!e�ir��#��3�i#>�#��(Sޛ҇��W�+�X2��"j��B�,�%AH+LUp�����;��(�������"TmY,��KC+^V;uul��Ի�n���w����Շ�����r_���C��\诫Sn�}��Z��Ǎ$7�?��y��g��!�{����vg�w�󋲎`H�@��t���c.s��������:�ё���K��*i�Mۙ{+h)��]��Ԫt��T��%��Z��6'�>�6�����;WQ��:/�*�~��+Bg@�i�kԊ�{�ڤvt^,쭃������ٽO/0�04˱/9���%H���
ѷ���jҧ=���$ݩ"q)��0����=q�#�(q��f�(��0B� 2/9��Z�@TYp,z~+�E�/8ܐC�(s���NE��:��ͬ:�`�N@4�v�p]��
Ԅ�%8��m���'�G�<�j����یa��#���h��W�� �z�x��3�S㽾��w�1!A�j����$��:���K�=�D����¹���3��,񉃕N:N�}��O
�d0�;.��Ka�B�C�"[R�o��B-J��'��o@�r,��o��s�7�Ô-Q�jt��/���c3�1��s#�j�{������ ��:�`Jl�r�A6�N1s}^W�o�*��䉣/�p)��@ruڃ��<T�?t��:��w�SO{�y��l��,�ʥ�j�L�}.J��k��/�������ڔ��b=8�{�� P��z�����c�X5������ݾx@��g)��KwԿ��ӷ'�"���θ
m������G������[�|��&�5Շ�c�<o�1������d�3�׼���;��ŉR/�_+i�y�3Q��V��솒�~������`0��UmZ^S�T-#f��9e�3zG�� [�A�ڷ�G���V���*lʆ�z&L�냶�v��t��ݫ�:�6>���6�D�:��d�xF4�C6>:v�"�1Z��j���@X|-�� %�~�7��H��&f��x���Z�K���(�]F]:�򌢺��w^�Z�;��%ݪXN��٪mT��-ۣ�h��.��
�r��1��:��I�Y�c�e5���v���$kb�}y�q�Ɖ1�v�L��r��p�|�s,on������0'uo"m���@���< O1��b}�(��b��Rg�Z鸡����S
���6B��q�Mȓ�<!O8A �DqJ�kyYW5v�3���ؚ��NQV��2;�(����>�ټ9�.yX0�]��cH�s?%NT��Ek�Q��`VH�چ,2No�/X6���j��>�,z�t�z}��.n��n�^�=����PJ������[��t���IP�@b�RA�R�r�6�ڍ>��{���>�����83NO����ʅ�7@T
�4*9[z_��Ul�Rɵ"�0e�{J�[󒜳fG�<��VZ�|ɱL����C��|�g�I�x�0�plt�>����}�K�Rp�"G�Ksw��3m���~~=9\vj^7����8\�z���	��5���=�CY��롵�G�<4�=G�.7bl�I(5��4��zK�.a���LD�\��K�F��_/�,��tuE�%�)4��Yĩ�����ߢߓ�!1	�ۿ׹�x����*����k�E����`h�Vq���OF3��u�]�Qec��>Q�����Y��߷U���3��#������C��R��im����u�s�YV?>0��p�>�,�
UVWap��=lk�Ya�^�������˨0��@x��¸�bd���35V)�Kv�Yg�یT[[�����}����᫘�4�l���[���8QKM+\�0y��fЮ.Kk��E�u����߆q����=��%tY���R�2W_�sw(p�ڸS.k���M�-q1
q��!g�]��ƫ�))%����nC/�[X>�������f��Ɯ�+ه����v�/ɔ���1�ٜE�Wo@2g@�y!>�F�J��9�ܒ�(�`��ݦ���������d��ۉ
��U�q<�p#v�}�Ǿl���{C+�n^�使g��!��aE�t��-YlbKπ��J��lz"GڦF��z{�&|@�W"���C/2p��a���(��#Mk�ōX��,�z�.�TT��3��X���Ԉ�}+4V�3�56A=��5���Z����QÙ���ܷf�IM5��c�f�6���T�k��!���zG�zb��xU+�{�=�✻D5ŉ�K�6��Ά�3�>7��K��m�-�T'���.��H\Gj��Ϗ^oØ��7&jj0�����D���4?��4��X����'x�ݲKr����5�bRZ����gX'�m32hӤ��e=�a�y3#�`��N�v2Þ_@�������H�%���x�2�s9~���:U�AF�x^����G�1����(<���&�O5ٌ����=2Pm
Mp��8`�����ec䀻ǟ2���)v�d���:�ׇ4h�1��X {���kI�����ɯz�t��
����<�%�����qf}�=�G���b����v��U!��g�9����Rcvd��R����V�]W�a���t�ap��xW���^ޖ���Rۉ��K�ځ�21x���&�~mcc��W.�bì{'�3��aϰ�飋�8<�/d�1��5��Z�V�`��$jg	Y0ה6�s����*ɟ�y�,��31��b��$��m����ǟ�bE�j��q-��Why۪�̖�e R�-a���2jPmɾ�z(�O���xp v�I��7�Ῑ��[�;g��Mm��Nr�<��Z�Hus_�H��uW�t��Q�(i�u�;	�ܽ,�b}8Y�D�k�Xmk	X�8+�X�b�*���*��GgM�"��Ŀ�@"-�u��L���GrckuI���侏�{IF�+Ǵ�5�1Qc��!�Б�	(O��� ���1Ο{�)�X�;�9�J"����w�zx���-r�n��?@��w��3~O�e��2�IE"�����+���t��zq��8�����X���~�����K�&��ʮ�C��<Gu9��}v��?���8Y�K�G����+���F5�}E6�'�R�qݪ����dЃ�W%�*Z�������Sg������|���?�X���c]Ϩ(m�m��˴��%]XFG�Ȳ/�r����������S
�XN#�����K�[�����I^Ώ�>�ȼ	�X���3T�N�����J�7�u�چ�u�"�l~������К �ǥ.�1G�o�u��=H��n`g^V��Ӑ���"na��Q���Ylٷo�Tį���VNz�i�۪U-���v/�_��fs�b��ɽ�h����ó����Jq��~��ki�;�l��7n8���ߗG�}f�}&}.��?�֨�9���6��	xB�I5��GlQ��+9^.O��j����5m$w.x��v�c��o��NЄ��r2�ﰪYF_~���^�X����A�������$�S��N��Z���o��}y� }��8���b��m��'*�q�Q�\"���)�vc��� ��ӑ'�'�p+��D���I+'�K2,�x�͘�!��	��|�\tM%���D�g6[J�V�ĎGl�����+Y|�ӓ�s9D� ���g�"���E��~��1tm�$��g�dw�m�ƪNtzEԧE����+��_�b0&��ei9�!��-v�)�D]z���X3�r��E�w`6�c��5�4!_�T���.����w�Y�����7���%�I��v�B-�÷?;�R_���	���ON8�1 (�B3l�������;�Z��F��2"w^3��ud�.�"��i�k��ꫪ�~��wY��!�y��������ޜ��M�9���R~��?�I7-�n�y�w��H˓g��[1	�?7��3��3��Q)������
��3��� �/���1���c��%4<F^�}��9��C����_!HS\��������;n�-m��hi�z�Afkğ(��R<��C��ɚY�ߓE��!����� ��R�����\�f�N�M��g�\!�8�O�q����ܫ��S�nL	i!���Y��P����٠��z��Lon��������)��1���1�c�H���|��o��H�v�Ԍ�~�)�\9��<�$�!�,��96n%8�������e� �Rz�Q#��.��l�kt�E\N�������?���Cey�{O@q��Ε&�����<q�����-����a��q��=�����LU {�ko��v����{�=9�ۗ��?�YRd�N-K�T����B:)x���p��o���E��"�%	fϟ���-�t���G�Q���Ѐ*�������S����*n��F���=��c�\��~��f�+��Ζ�Yl���>J����*8�:&8�6��ot������Y������o��V(pRA��m%��W�`HN��J2��@�KU='y��i��9��;I/�~y��w��z���XF��k�u5���_�K�����W_=��{G;>� v�@����9]�cC7q��`��0���x��Q��&*ܪ������jJ��{�[����*���8/�Bf��=���-��`�\I,��Y�I|�A����M�c����V�3�Ԁ���2V���jR���Ԑ����J	��G���)y 0:�߃��:�}#�=پ������qb��]�a�t��qC�\L����uK����iX��8��z��/�[`���YeҺ����Ƭ��%��Z�M��H佧�t[���[�#��v���y���%�Ij�r��u�/M���8������������p���l��[q�~�v�{@O}\'����ճ1.��o��^q9gPE�W� 7QO֤0�Q<ǬN������L� �\!>��٤Dѥ�F����5�
�_�rv��/�uk�p���J��=�{ �annȝ�<�ȳ���?~�Pq�s�4��U�Y_��ߔ���ڠ�t�[_Y=�?������	���4��`�oF�>Q�Ŋ�I��Q��Ʒ=�o�{Ή˱�����+r���滩"���%�?:O�O���G M������7-ң�x.I�/7���\�J3M*=�dN��u1��s\ j),��Z.���N��SJ�s�z�ۭ�4#jc�U�Q9����a�|dh��+<��w`�2���S�;�6��՗~Η;O�s�}#��v�ɑu��Y��āB�o�j�&�"-������9�P��`L���r���#)N�p?���W<�{�ͲD�*9�醁��6P�V�IY��vڶ*��ǡA�3 zv�7&vT�H�S�%�.jvO�{�y��P:ac��9/�e�M���p����#��g����ob� bȂ�[�٬#��S�;O�k�BkQh��*��s[ �I��.ɓ	(���*)�A�H7'Z�_� �k����0�a��p�ף�4ˊ����@$�*���7����� `i_���ɕo��4�1��4X̓���rjH��>��9K��s�`'����f~�� ��$���G����tN���w�a'/"Ia8��S����V�!�iO��n���:�,wk*.��el�	�� �7JHhի�ʬ������e#Cb�)~�3e^`����O��ä���%qI�)��[%���R� <��~@\���u�&��`f+ň65e+�D��-͊9���e[�5���b�Uc@^��4Ǽ׈�jc�Mv��;H�����͵�J��х�^3�V����Ϩ� �K㮕{����mt�0/{/�0~Q����JvY����}u��J��� �Z�p���«�ƻ
\�jM��u�@����������H)�pK��Y��l��~X��{���٩��n������@qEBe��2_#�Q贄��/����"`;	1��nޜ��[� ��[Xi���v���ѧ �C`�����������2A���e�*����і��ٶ�Py\1�
'H�ֶ�6���� X����P��qc�->]�Ȫ��T�Ũ���r ��<.(|�M��|�s���w7��fO���=���#�	v���~�!O�qZ3!M� 2�hR�����c�E	�V���%���$�TL���h�̤u��	"�
$&c�;�$�~R��d��)v⡢{�;�Z�@����������:K2����EE��W�P�B��b������=0�km�����S�.^P��fr)}�R�&H�ʤ�����~D.��q%J�^�5���^��щE���K6ɞpqȘy�T,�-������/��T�'O�_���xs����-����\��b.�5iƙ��b\\*
�m�h������v�d}+��vZ�e�#d��䢻��
�){��L��:�-b�l��߿����Lb�D�!z�l�R~"���{�������<��{�/Y�ɶ�hR��P�{w��A�H�Cr�n)`�RW�{�eRUYS~9q���aK�O�S@��1��.�ր��Y
�hz��9�;�C���#�F�� ^3|3d��!U��pY(_�;|��sqN�\������
t�)���F��]�_��I�X��4|����Ů���Cy�.�~%h�O�Y����7:�����k5}�(�.$��� ��8�iQQyAo���`)�M~����r�(s���{Cˬ�|P%�~_(U��*k�.�9�[<�<?���7�a��;1��b/z���?
Z�Ī��{�  �k����k�ju'����ٻ!�"�5S:;	R��[�-b����������_	'��S1���.\��%�;>�`c�+�`fg-PX�����G9{0P�E����͖�Ǝ���+$�>�_����G�pe-л���g�	��{�(9���tE�UbF�
Y�?tP�jo��C���E*oG�^��1C<)�@��0�� �W2%�����dj ������E�"=2�@WA�B� �7���.��GA�wTO|�:���Y�F�5b�3��#7�A�� �Kl�66�C���\�4Qt,�����ц��#��.0x=�u�4H�/-W��^�R�5ۢ��~�z��������&qw�s�(����?�s,�we>�=ê>֤n��P�C_��Zv��u�Y��۟���v�oVt��V�};}�Պ�	����I�=�<=��.&�`,x-��m�}Ԉ_�.��}�L~Q�2�(j�tD�+\����.���52N~��?Pm���׃�d��X���Wo[EAޮ%J*r�Ow&��sV<����f���a��PWR@,"T��vtŢ��z���G?�dU�q`ͅ��U���ҵ�I'G>�JȼF�N�n����d�W&����n�xD�K�C�O��qw?)*�BI^�ɍ]
�?�g�-@�`9�v�ۍ������:Kwn���W�A<9f�1w����>g��x��H�8{;U�}X�@���E�/>���o����V�k���DU�Ug"�%K�+�}]ED���U�~W���B�j-g�Ɒ��*B�t���3�"F��8���D����կ�|? u>��R[�֐��?iq��`*Ef�V��74�-����w�C��m�\�Ĝ(@�|�W�!;��="��p�G(�*��6��]�	�����~����W,��U��P�i�Y���|���������A�6�au"�DI<��\�3t1?�����}P�,���� l�2S�F\+�`��; \��ۀ��T�EѼ����ΩL}���I�z�7(<������D���r$FP��v�&yn+$�'�D�C����f����ީ&7����b�!7)tX�^�⪘�[�(��R��9_�\6ʩ6�%\��ץ�|�i�ƈc�$ζ(TL��Y?�O�s��;���XMkD�s4m�B{B���Kޞ�v�*�Юj���S�k����f1��Wu6wbx����;6�M�G"�T��6������l~	�=�t���D��6VӴ���Tά�_N�% �ݾVRb���N+r�t�I��u�da�wvy��|x}0.w�����=z[�!���a!{��? ����BeB�	���!�B�ƫ�Z�V#��j� ?�|�� �P��$Ue=��ό©ފ���N�<6'��qϯ:��,Yʒ��b���` �<i��
����p�D}���/E�� ^�f@�?�}A-��c�����z�9l���R�f�`Vc;9�E�G�k]��p���R�J��`@��.�쬑Ju��ȁm�9.�9I=z*Q�f5�W�z�5M�I.u�ZE ���M�Q;�.�k_����kQ���U�l1�H8;�;��#�)����#�@{���f���� �9Xz���.����֘��>��3�����e�K곁�1�s�8o�sY���7�r�E+�$��_��ӯ��ѧ������z3� ����ٲ��P//��R�����<u���H����7���e�v��|B�
�޲e|t�A��y��4�K��3�$��7(��;��n{ '4�_*�x8Pùo.�V�p�w7i@D��"t���,�BW�5g���.�w|����J�׍7D���R.`g7<`��]7�rF�B�ׁ�J�-��EV�U;��h-#u\����p/þ%��ZpH���y q)��e���qk}y�GO� �u]L��߱_\ء��Yd�<n�i����
lO�2&�b�)���A4������f��W��� �w�X!��4��rY��@n�1!�AW޶E�cE\�S\��e���A�N���Sk?�J*:�]��4��%vn��z�ŷ5W� �\�z�
sݗvC����t�L|�@ L�k��L��.��o��s)j�l�%:�46��zp+d嵼�Ţ�K(o�H�L�V�z&���[�Tǉ9
xѨ*���]�ʷhji�g��"����.@u�NYR��^lK��x�xlG�vVz1.no�cI�hE��v��\dYeY;������$���y��g�(�j���tU49g���*fg����q��gQ��C�s5�����}|ڴ�]�B��l�����x��ܕ�T��CeOY;`�̊��`����Hz�շ���\��ό�Ծ�� �!�.�H����?\<O�lM3bw�d]�<����Evw��74F$pj�w`� �M;��!l#��;E�k�U��>۾��R.������J�~���X�Z�U~~Z'��BwxN�iÝJ��l����V�)�ۯ�'2��'�q���\�{:��ZQ5[����s�M�^2$�k3]W���ɋ9���𼒵Ν�9Z�''�	*��K.�#ͻk8��,��t8���D���F�m�z���ƽ89މf�u	)�}/,*7 Ҭ.�6�:g}��w��S�ή{�А�x,���f����*�B��/�w���ZZR�v>�3�:*#T�u��;xK1�"�k��M�H�wZ�i����0�⤃FoP��p#3�
��|�L���:�l��%[�Ky%�냘��e��O�i귇�O�Dht�P�/~�3l��B.��RU.��~�řk�z��f֔Tu� w����<{����>��1z�g:ŋ�x[R�<4C����b`(8s:�H�;�@������ypG��5��X�6���k�1�|��k������m35�1|�e��˯Ky�ݍ6�`w��{td6o�'�}�fB�^R��Q,~�k��6�H)��l��?����v�A��*��g�s�b78���f��Љ*�m�Vժ'�����SZ��^S��WD�ƛ+WT�`��A@ ���6��u��w�M~л��a_�jpB�Y�� �ݏe��Z�0E^��7�@#کU�ϣ��ҿ_��*����_$'һ�r��}�~��M^P�C
^���P���"���J��\�^�૓e�+��B�f!�u�ޗ�eUt�M�7N�&�@�.�s�v�уD�{�[��ocB��#Î������c�2�q�ȃJ+d|]�����9�+wb����c��� ���M������Գ���sg�Qr,~}Sе/�g�+P�w�f�8���-�V��W\���~��J������n1�;2��\Y���T�+�t=�u5{iuX�����$s�%'��e2�q����۷*%��������}[2��M�Y�ڛ-�֓���0�w'�hR���,<��1ԋ ]2G7�<������F�������}֩w'	�����z���;i�qR.+���e~q�в͸c#�f@��Z�eq��f۱�+�������B
|ܠ�{�c�U��.\j�c���Ä��\��k6nQt�k#�ً?Fn�~��o���̘��^q�}��� �'��p�^�W+���4 ���h��͝!و
XNV(Z��蓟��~{'�'��ҷ,�v�"D�+Oغ��]��-t�D_R~�q�����Ph��N^r�_��-e�J�Uڢ��r�V�f����'�z#���7�@g_5��� XhKyHQϣB�9�Q~����i^�c�b=�J<>�p3�y��>����~ex�Eb|�+�_>���p����%@��?����~Qww9��\���3�� ��Vire틑���$ε�� ��3<��Ι�k��00�}�Y�]����[��4-\�
[��j���X��
1Vo�	�_�*�9F@���4�I��p���i�x���*5��g��Y�k��蝁o���5B�j�{�`�F����j���MjGE'WH�6+:��CO�F���`�&׊v�GU��@�������@��tiJ}�~o��IoIB^��Mp��f+�C>�3��ͨ!���J�h�m���K�cǑz����3��4s�����lE�Hu�f�md <�\A'�L��D����{w^M���g��-�P�֗	�ׁͣ��Ђ��ǂ���.5!~*Ë�'պ����q}�
 �7u�`E�M^�#:�n*��G��2�m��~R`5?ЫX�(�5��X�<����c�E�.���t1�&��,�d�`���k3��6�*����P��W=?�ƍ� KrZ�ؿ�����ؒ��I�r�q��»D���J�tM�b�<�j�mp0�~>�vXΫK��8aH�m�z$UN��~�{&um�2��Cr���1O��6pj����X"��o�ޯ,~R�;e� �l� ұ+���t�⢸�Y�EE��0es�qYVHw���L�n�KT*u���pԠ�:�&@�7&u!t���$��\[��Awm��_ܺ'�Py@ɸ����� �1��f���e]��_�(kR���n���FM����y`�~͛��}����|�F���޵��2��k�,�@>I�"��B�ǂk�#F�*)�bT�A{	��M�%�t���4�(��mG�-/��Jٗ}����D�wa���W�`�Uxb* �������*8w2ݟM�{����l^����$f�933����E�z��O�I��
j� ���5[6����+'���$�x�r�����qtzkmc�?�DuCf�&F^�sO�rk�s'O����oG�i_$��|��W��v=��遅�S3�FZ�9�d1!����0�U^(�"�UA�H>eS�H���<�tQL�|$KeZ#�T��e}M��J������i�I�x�C�cQ������P��!O��J2;�VSF�ٱ��ݜ��"q�[����� ��7~���4�نϷ}�O]���)
a�q�f�{6�Q<���y�����g��S�FnI����$4�	B�[nA���Ěl?�&�2S/J$�8�]�v��v��V���p �\T1���ў�4*:�vu2����0 F� ��Tp,��[S��`6o����buG�ؔ���$(Q�+l�*���M��Tu̶�G���'���k��*�0i�`%�F��#�D�x�0�gia�噐�֗+[�1��ئ���+�4�r�%ǥ*��	���_ȫ7&�5P��J��A1*~���I3e5�D�g�����lUߊ��dWζ����$������+��7��/m����r�e�����sy�m��]/�70�69e��t�O�9c��B�R�����jچ��mZ�P�/�o���Km+O�4Z���|*&c5�w�Z(��Uږ���<~�r��fN�p���`0����U�{��v�i���c������>���_!OZ{�(
I�Z]cQ���5���-v�:�����g�W���
�a�U�{�Nw�{^��e��aMsJ�s����ӊu���c�~\s�yJ�g���&����K�2�&�zEH5):RǷH��K^�>�P�����~B}\���D� �� �����7�N��}_�oo}��$��V�+JJ���z7i;��I��j��-"x~�|-���HgbnvT-ǲ��(dK{�F��o?{)@QL��\�]�]9H��'mz�+sk8�j�%qE��Ee`���K�RڔF�5g��(mu퇹F��i�-���v�o�yq��-AF�r�3s�E��9ɪek��g�SY�,s[#�*�����l4ٺ_�$N�4�c)K��f�CF�/��"��
�6�4�W��+��(<:����u�&��I]�Ď��0k�}$=���/����C-�4�7��k�P���`8��8"E���)�@�qY/c��>�{A,?���f���4"dǼ�o�������l��G�������?`F��^�Zyum�O4ױf�'�,����~�wCUG�n�Z�K��K�~��+�YhQx���D�8#|Z����cLK�����o�K����j�]6Z�F�S�G��V�c֝Ȥ�WQ�'24Q��rKԷ$Mθ���╗�C�jS؋âق����v���cv�~+�0�}v�gE;��t9g=��is����<�)����2`�fy\����|nU<��_H��	:�\H Z(Y�$a}�!�c�0�Q-E����W�$�:��`AE�+q
�|���:*�{sb��Zxf�Rr��/\d�
���7E)��1�@���.T�Wa#3qp��&8�������E�&�%P�b}i�5����rη�N�	����h��3��>j�^�\��wB܅�S=���W$n=��1;�r�w�v���M=��e�:���Ҳ}u�Tq�_�F�_Sj��dٽ�Y �?J�'��=�1D�}��{f�z��"�������k�f��s�ר魵1�j�j�� ��P59��m�D:�3�@���q8N�w�� WA�?@��	�'0=~���މ�|ڭ)���
��v=�@Y̖����Nn�ƱꐑZ?#P\��	�jj@�'*�ݑ6�غnW���Z-D��	$�������]��݋�Cr#�T�{؃�߮�yX�y/�a~���A����)ٸ��3#����-�a'԰,�)���1�K�n��r��4Ɋ�N��@�'n���b�E�aU�������5�"&R3�H�z�yᩎ�V�soO��<��8��>W���$�q�pn�룔�����"&0J%�˱Y�����>�Qq�r�.3������nD��`��$+M�7#���"3�B�xV���HbǞU������|��_�yա>�c�@h�����_Y}�ݻ�A�]_���H���Uh*`wN��:z���롃<��}\�f|���ve������C�7&����_����EU��xCС�J�Lm���+���`�/�
��2����k6[��;�v��.���{�#��֪�h��K�Jճ�[l��u���[�2/|�9�^��/��9]�W�+@變 &&���o�ĖU�h�Cј�5����l���1j��W��A*o�'�w��T���")&]O ��bm����[_H"����b����lq�ܕ�J��@�Ow3p/l`�!'��aW�����XX����x'h������?�Y$�X��ɫ����v��%�y�z�Ԕ���D�a�e=��4wW���O�e<�]/�h�|���2ooƿiZ:>�m���pN�+c��-/V�	6
^���͵l#jA ���$�z�8")�+�i�r1Z-����
�cB�&a�6��fu�߼<ԴUO����]�KO�4';�&�,��\r��'J!*_����Ư>�ne���MV!�D�*�XH2�vo�V����a������M-G��:��.>�lH��z��o�[�X��=���c��ܧ��M��]P9_p5?m9&<�(�jv�J�҈P<���㳝oqk[/�nLte���|�k���i��f�jI��6�X�Ja�gw������͐ �ӏ+A��U��<V�Pg�XLupO~'Dc9\�k{X�2m����(Oyq�,��6�7Dbk��험 �b��~�$v�Q�)�S��+��PA$�	��Y ����&�Α�oOl��7d�_̩�f�;�I���G;n�}G�ˏk#���W��A¸���:�A�c,�`�����;! ��F��G�}}��h���A��î�Q�\�B�i���Ogf����vn���렟�t�����M��e}���F�k�}�8����ҝ�]�iAZ�{t#���������������b��8��y}o�v��wg�tj%�{�_���O��3._i�L�[���Q&��[Gz�be�MX�/3y�P�s��e����;%��7�@��fIs�,���>_h)�:ʃcĐS����>�Y��l��c��nlJ��D��� ��UYIw�̂�����L�C$�v- �ȳ��"�2e#3��4%�IwQq�� 3yX��Z��D�$g����p��.������n1o�z]ht����n����/�7&cN����Y��%q��2��9���r׶B�	e�9@��E8�(O�+��0���K����m��#�m�����l������S�X�z���q/�
�:�4�j���H|����I�Ϲǖ��̭7��E�hTr,�PZ�I�@�͆�2�q�G`��߮�[f�������:�f)(?�������P��t4]d��p0Xv�ѣ�Y�Ө]�9of,i�٣1��ʾF�/0t�^J��w+�m�1�ʬ���,����Ԫ�Ȳ��=ʕu}.�ؼ��>ڐ�t`�"%����X��X�Y+����$2,�2�`O�thN���-Y�,o-���_�	8����l3]���*��CQ�%L��H::����ͥ}Y�Շ����	|'�����kq��C�pW��s�����eJ���o�@0"	�g�cɫ����._L҃3���}��,,,�����v���R�g�\���=�zL��5ɲIΥ���gW˒�VR<S�g�Օ{��o�s.�b��<M)F���e$̭�c�hЫC	��u1�<N�0�G��!�M����N>�i8i0[ϨG��j),^9)L֙����^`���Ե
'ݏ�F�C9��mKf�i����B�/�[�;f��_�hC3c2�.��tC��ǝ�4�3������0�\[�ˍ�/O}��e�����;�.��Z^�v�u����4��G�AY��n�7-l��=c�n�T�Dc6�w�Xߋ�~���@���m��@��$r�|��>*�Q�2u��ҳ���(�9�#�?��-g�I�z�C�2b�C�~91��-��k��n]{�x������{9lT�Ջ�ϐ���r���Hð6QS��g'�����ٺ�>��U/�$�;�J�!�ɘ��}󄞫�{9��w���p�<7��-���a��!��R���Jd��I�a����<e� �AK��!�R�y��k��e��#�Ͼ��sT��u�p�	�=�iz�:�#�s̸k��&)R9�^}c�J������;XyX��;��Wa�#͸U�V�u+z��G����| �3�j$_B��Ջ�@�:,v��X��Q/��@��Eފ��L��)Ί^��RF3�U�����Og����lg�'R��j�A�mj*×y��S�d���@�:�^=�'�ٷ1V�⒕a���E�����ҍ��;.[���������7'խ]��;N�ۚ�<*F�p~�}YHd���u�@:--g��;���������扆�i��Z)��#;��{?����>�%��4����<L ?�di�ޭ�	؁ڌԧ	�����U�Q�^}~6�'���{ڜ��	|����y�d��A�f�6+�\O&n���ܾ�:��p�}[=ֽy��b-�&9�Q�0ǅ�>+^g�6��\�yy	S�XB�����nN~S/*���D���O����ox���q� ��^�*��Oٽ=Is�M�>��4����.]x��]��YRY��I*=M��G������z�\�e&K?u���
�/^[W�n����b�k}군�*���R�c���NI��&o����C�וY��к8���a�� ^ן�C�$��c��`ħ��$�ٚ����.1L�v ��c��^���:�����lh��m����̛�^��Jǅ8) *��ᒅ����^�|�]�{!�v;·��Ƙ�?��g�����%'h���v�A��� ��	}9L�hu�@#�ƿ٤���>��f�\����w6�n�F_!���	�Sܸ'��<TǮ���Dߣ�׉�rp�қ����^���ޡڴӌ�#>����u�I�D��~������S֎����N6����jl !يB��e�-��{��럃v�I�C$*�����
�m}T��Q�ә~����MEsɔ�;zn������٤Aw�âe�ңu�1r�C'������}�XƇ~�yvGx'��w~�%�Ҵ��8�V�;�|��CGq�c�x��2���/��`�׋��{i�p9��Źn��W�t����N,�k�#�}�R�=i�o�R��p�7��̖��k����m�-��5q��ҭO ��;���{s�ýF|(���洭N-�����l�_���!��
���e�W����N�`�v��X6���G24�6]3�R%UP�
�3�O|k�*4wWP�H��C��4`7��$����OX71	���z��.I����uw媵��W�	�����"L5sn���H:>HNZ;��.Y[��:s��NJw����v��f"����߯ŵ��������׫�>���� 4�~[��;Deo���>�Ʒ$tAHȢ�E�[���W]r�� ݀.���Js9mfˬ#��
)f��HoD�57Hgz�� ���o��D��g��z�*�H ������6|	�x��
=�U�K���olQNq��Yϥe���b����̄���7����Q�'-IE�f��_���Q�Ѽ����ϛ���Q��ዞ�wS�~�{���Պ�u=�=R�<�چ��og�B�@_g�"Ӧ:�u.*dg?ŝ<d[s�d V�E��J8nx�4�,aoڿ�z;�Ǥ!<J�'��A۽�0��n���
��$5�Ook��1��&Һ��<O(Z���Yt�i}�5H���t����-OV^�w\|ymF�a�e��4&�F�~�v���| iV�8*�Le�*�v�5<X�V���-`b�͓u�����Kp��E�l�v/��CQ�ٮ��L���L�}|smB90IS:�x��$�ɑo�y$lwU���^��&j�q�$|ȃ�f�N{�L�uJ��ޱ(�3ˀe�$�ck�&ˑ�ٖδqh^�"d$|��4,Lm�#��b�wJ������p+~�.
>~���d�?�Ŵպ���A�S	��#4�r\�3�ZNA�|=q;��&��h��{�]{C��i\|���ݐ}%�αx
���n���lC�0֊��e�س�����T���H�,��
1�Y����e�c�گ#��u,_W�67����'��@����+����-��%^��eF?�*C@��ɪF�3��*T�.��φ٦v3�[�?p�[њ�Æ����^��2gDG�.��c$X,�ƅ��:5�k仇޹l��{�%�3���i�>8�$�����Dv��B���VJPh�'�S(���*xJPϖ�k��I����h��|�OV�"��L2ۊv�*�M{�4��7A`W���5��k@H`>}486�D���M�	�GIJm��~"k�u6����a���ay��?)�����
2�pg~��>�?p���,v�-$��2>y�MBA����R`z�P�q�h^�/.����<)������|^qxr�y����drR��i���f(�~/x�V?%��=�W*��:VL��@����N�d8A���L#��χr)�pyvM`��o.�rf�0�������Ҕ f�����H���$��+�"T=��.,�Zd���k)�%J�Ǖ
�B�(�ӪPO-�\n̏����CRs8�_ɟ��2�?n7�&�Y�Vm-��ϣ2V��(h��P�
s�<�����}{��%o��(�%��'V��Se���d��@�����8���*U(	�c%�^z�ya��2�^Y> �j�u�jѧ�$����ruF�5�������<Z"U��,[~���o0�1ʪl<�?�e>��8�m�NO+��R<~�d^�I���~�����^=��Sȯ�� �s�]oSU��Տ�q^�m��(!� 8sNN�e���ܜB���ܳ���S
��c-a'wF	���+���<0��ZE*O�z,���8�-�0u���f3C�*;x_��'�8��WQ�z�����U�i7oqv�[��,�է�{L�ܡ���DrH�#?&���Ա����D�u�!�,3�r̳�"!�SkF$�g��"E�DV0je���]T�_ĐX�
~�ڢxd��6U���HIg�O����G*5O*'	-���gl�Eth ^�K�����
�g���8 �˖�5|�"]��9�p��X�[�H���L�n�-[�:�+�ӷ�^�_rC��F5� ���^��G7�W,8�63��MBY5�7S�<�Q�A*��TO(Գ%by����粭v�'�a+���>ߏ}�}����ɳ
N#A�O�Y��'g��#!m�%
ܑ���`�TB� f���^�4�W�_�O���2���ZIe�2�[?�����'�(�DX�!��G�k�8;wda������]u[�_Zb����̤D�:��X(�Q�kcQhS�~����3���O0��pwDXٲ�[ ���{b�G	�6�3 9b�e�#�������ݯeM�ۼM�K �O���x�D@��J�B���J@��dm��C�X����Yƌ�O��~�ڽ��+�u���0 '�1�U���{s�SA�����n��;���>?�L0�%������Is�$t�˾Ok�� �ڮ�*$Z'�?���ݮ���.����l��P�T�͓\�Y������W,�Pc.w8���*Ux~��ڱ��dd�Rd8�_�=��P�-#����WP��H��G�ث�y���L6�!��de��|8���9���G�����:^w)�\�?,L���kV� ���PQ>�c���>d�	eu���}[ZB=͛�]}��֭
��M�	"�<mXB �����O�f u{���
��6�[衮U�7�n��/d����	��*�8����Y�)nw��)ۀ�ٝϵ�>+��~��߰v�a�|ʞ���������"����|�ha�S���?\���}��~�<zٗd��{s>�U^�E��3�s ����,{�#_\8��dk]go܄��a����3#���e�a�<�����}�d��Ϭt�	�P����0�W��.�qe*��.�J��Z�ˆ�枣�i���	�����M}3�@����B�48���{S�vl�.�
Kov��-�':��蜁����"�8���zv+h�6-4@�߰����1:_ŀ�
�nqü�f �}V:�q���]r��:�쁒P Ժ��Y3?�]@��ӵA>5�mm����]+��W��!����|��W�n�ܔ7����#PK:6Q��/B^��kz����S	,3�f����T��l���i��="[��-��4�:L&�rb;��$ᜢE\V�n�'��/�0�!�r	��ob�zÓ����g}���/��Q�Q�RcovWG����a����@�Up[=Zê��
��u�A�i��6�X�C��x{?i�$�D�s���,u���6�huZ�
9�����5Ϗ	ӑ�E|��چ1~g�st�ˆ���!����a/���������L�/���.	R�E��*ݒ^Rd=Ѽ~�ghma����,91t;��\�>N~�n�YA���&il�,n�v���R��ϿnT�w�Y<�/�������?6��5��S�d���"��1���4�I�8�S�E-�p�SyT���H�Z��W���(��ۙ,��7כ�֙��.��:N��kC��C�p�'2M�T"�}ԁ�"e5�]�;&�MiB��.o��I9饽�,���&m;�g]G�t{C8����[w}$^�k���侰z�(�������X�`�C��`��j�ʏ ��O��VJ6�@s���M6i�3�5��"z�=���9�e�Z�P���r���P��]�+׊>z���c=P쏛��c�})u�������C&5R�ڼV�PQ�N�����3ԉ����6����G2(�l&�s���������[�l���w��2�[��H+؄�A�U��]���;+vU��)bGy�����ޜ���:���� ��4�ä>�u?ڞ����-���:����ޫ�k{퉺W	W����{�.�ϓQ�U�>�D�à�Qq�j����g��nx_��ci�ݙ�I?���`���pF� �������犓U�19U�Zӽ�uJz����[H�u���3���N�88���!&�ůr�p���d Xz��!m�j�p�]���r�|~sSwvX3�x���
n�tJ�跖��x�t�82�=zE|�%(�@�O��d����WoR}�K�݀�������A-ϔ���$R��9T�z�B�rG�0_j'�pa"�倉�7ȹD�@XO��.K�5�����~�pTAj�'�_�s�~��A�}Y� mh_�/Ɍ6 �=h�b%	Ɇk���E��q'�il�}T"Y�p{�k��t����;m�>M�z�'�-�Z&�f?u';<�M+���<1�q�����
��4���q�m���i��WK����B
�l�ԑe1�w(@jZ���9���ξ9�\2���\�FN?��
܊������?��`�A	�i��ځ����,���Uu�Oy��ql����)Y4�wK����=��^E:�1�>P����x8?ZX5�^���4��W8�U��4�ډ���H�$?�&���S�����9`�ON��=�p�݊ ��ޭ��`�����콩��������Z<��&2�g7_
^7�ߕ�>��"�^t`�x/e?��t�q���� �x".*y�C{�Z퍪KpB�Ex�C0��F��3|pz��R�=T$��uvZ�U�������} w�ҟ�����0�u��a��~��<��]�A�9��{���Yk���V����A��*#���%lʤ���B���6�]�!�:-�X �̇t�&P������~��#T�r��$x;�D��	��5������n'￿�&��V���$D��	CMp����b�`����^Ӣva2w�]P%�S�wQ�|A�&A^h�V-�M^ ��B������?���qLҕoV�������)�c�*��������D�g��n��l�0I�0�$�����E���tA��7o�n's��j7Og��A�Uo�&I�Z&�o�Ӕ��%� �e>q^����wr�m��c��/k#ݨ�5Je��٣�'|-A���
��60��` ��|�b�H''�9�|T���n��σ�/xCV�%�({�����\���-Ҫ�T5DՇ��ն�'�f�������=��a�L��?��RU-P�*r��n�+4�zQ:�M���x�>�>�����D�aI�ߗ���N�O��㾆��?�7�:-�9�::�L\��p�7�ֺ����X�u?b����p��O/;y$gkW=Y�K���#���"G[x0~,
�<����S}y ʬ��Ϥ��+_w��8f��2�L��AKj�9��<�B|v`�P�n���.y%pCT5�O<NS}��@�|!ǘf�z��G��G-:��la�?Z���r:�9z���!��4F�벬=u7˴���gemOX�8ǧ��בM�=�z�Z���=Aϣ%{�J֮�Q?43��Z�eF�`���mE��D�R9���[�p�6�q�b9�7��ma[��o�ǚ�׈q�ű(�]1���C�8.��/�u�d�
0��S�����͗����x��x�Z�����<um��w�����Ȭ�-�C3=Mi��cW�Wp�8�CF�Ҝ��[��φ:�����_\dTV��?-;}��{@�������0%㝦hɲ�[2 ��#��6��=�C���X4���^N1�pc=]���>
�C�����{�6�k�8�vI�5O,�1S�B�~��0�#�5�F�Fg]M���R�{�h�8K��H���ГӶW�c�7ڷ�����߮��2��3�D���l���3ƌ�bn��ܟv���aܽ�����a����`�z��dE�x����U
ɽ����1��u^��mo���"��܏��-���9C�ij��(��-�"�K=�ҽ���y�R5N_(vvi�*��j¯uA�k��h[{_�g���J�w�g���>B>'���N:��`�*�zR�D��4m�[w��¦߬����<\�eެ��rst����?"�������1��o�_�K�DT�4��a}h�`H�O��6���Nf��u �%�ߕܵ(����f�	���J��L�q�nzq?Bu����uڻT�6~���{D8�#۽�&��%^&��p�VX��<8��0IcN�Cc��B7��Kk������2�lr� C'ym.k�(S�B�%����E�Ԗ��l��h��R٤��ș��p�u�]�n��<��<j�ҊU�N{�^-�5T���Ź*�P���w�]G�������z�7�5;�~��sia{Q'_U��~q\y1����K�-��2���D�o�p�?������n]-����W1��@RX�wS��1ɀ�T��x�f\D8��.s�&$߬ )��ȓ��.k�aK֩�hё{n����h��bN���oMr܇���,�,�XNCT�p_�k}����Uɬʡ�k�̊��L"�ח�>�i�4f�����l����<[���e��w)�+|��s6#/Uq���V:������%���83~f%,[Q��R<��ې�&	9��T�Ƣ�%] L9�秌VMU�.P���>��,�Ζ��d�WC5G�7�Zţ
mli�waM"E�m��8˹8���'yf7g��6ZP Gxt�z?�ְ��y�2O��kko�io��4 f�}S�V81A��^�����:��4���yP�|�HA4^�����'n����7H[�E���O�Qju�Qg�r��齱;^��z��˞ɷXj"z|zq|w�I�V��z��CB~�節�;+I��96�b��J#����q�F&��eY�q��h���}�'4g�2����礣<7H㫳~UI�+~�*��m�쎗iq{h��)��Gn
��]"�!����Ԧy�o<��ӕ�ۣO4\&3_�
�VE����*�����>2ߢ����.����0Re�@�y��F��ۑ❭��ܣ�s��\��76Hk����¨j�P�6,s�h1�3{(\�n6�v^�k��}��A杓|"�"��]�AI�	���l͗^ͼP���M��C���p"-]�D����F�)%��8B6��!�%��]Ϝ��8����E�;���j�m�2MI�/���{��,��B�Ƙ�&��)�(�^ΚK^^Y��_�#,us{|�]4�|��)U<� �Kj~%��IF��4�t [��2��VE���(��Yv��~�|��u�I-ipr��ԧ�w6�Y#�[qbfjyr�����в�+*�#*QǢߺn�\t!ץ��u��/��W`!�l�n?�ʬ�GÁ�����k����ZuA�ʳ��@Ȟ�k��K�\F�ڐ�|d{�Ⱦ��3|P�2Z��YqP=#SZ��Gg�{�����_��҄JB+����=�n8靧V�5�v��Lu9󖿑���� ���!���gWw�l��abPS*����k����_2�6���Tg��Ɛ��q��̱�J�ş�Uݓ�{�h��Mx7��4΋{i�fFz�ǚ�1lh�S3��Y��e�A���=U�E-��Y�����
Sj��;��0�cCǷ��kD��<UB���{{W�\���Z��;�I��r}P�grʊV���8�k��6N���wי���\��׋��wf�����\~dK�]�5V����|�_�G:NW��B{��?��6��d��ڊ�.�槚�Q�������v�䈪�s���B�O ��gz�'���*=}կ�!���m��8?;D�7<��>�']!�����U?5.OQR`��>�_L�>3�R����
.�o񘑘�=B�WE/�x�:���v���7^�<�M�����@�u�-B:��K����A^��ff���, mx~��ۿ�x��������C������
�o�# �e����K
؂�%c_�Y1�+3w�	��B�&go�J�gLo�6)�`gC������a'b���x�E{�?]5��3�Y�QRp�����J������a0r�����xPpyg��dsy�.G�^�?�F˅��S�?� ��|ZN����z���U4�p���F���'����o[)�����p� �l��j�;�+���P	�q��+p����߇I(Ar��%0��YH�mQÌ��T��ΨㆸΨ�o����;���Q�� ����r2 `�r�c�����q����P�K�s�I����V�ݘ�|��;o�kh��K�9��x��񰯦���s�_现���n�C�DO���B���ԟ�^S!O�n�N̰ho�O��6�I����h�\f�;,Gw����B���>�.���2_6��UHӬ��.ֹ���Omi�����̾`z�ed�8)��]�l;s��Q���3 �.(�����]z�:��@ݝ�������
�q"���[Z���fo,����/��.E.z�=ˁw�7��S�7���-����j�����DQ��1���iIkW�L�4�P�sp�5˩��"/��Uv����o��\�99��,�������i��FK�Wx#�9�AGVV.(W/�+7ڻ��l%T�	�(��NBL�C��xЋ�j��yL\�p[Uj��.F!��?��jʢi�^�#��*�$� v����'ۛYN�VF���~����4Btx/v��J��������r'�d3�طb���e�dK%��Cw��Y��2�<LNY��b3�4��֒U���S�*��g�-,�Fi@#��l��%����JԷ�_��Uգ���)�d�wr*�5�5I.*�p-ӓ��Ǭ��Σ	��R�]�I]?���MW�ؗ�,�ɬc
C7c�����&�	X���l�u��k��6��|<{�^��d"RItf�-�X;i����'��'6���G{xꊲ��p����"�[�����N,�� �]���O��
��q�z~�ÜN'o�/5ԩ���Ǘ��P�%�{��/���X�b�T><�/�~��=s �5�c!�B�O�L��f�aS������`+x���vf�<��[98������GW���6Nm$�.�-<�Pe�V485�W�o��(�<?=w�|�h߱��œ,�c?����|2;fｋ!��)F�A�N����	u�O�j��A����'Qi��i1�ߦ�%�v���A��"?�	`�JOx��ҏbQ���g���2�"�u�f'�m*���2�)k���6f�H�/܉@����ԛ�ܻ�ʌ
K޺���S?~b��n��f���;4�H��o%/��*���k�QT��/u���v3���p����r]�a9�1�cB�]���zu��	ޫIF�©#2�(���R���r�)Ԗͷ��:��}��cy���Y�)q(+��+��Y���[dȴ%�,Z�~���u���[���R4
D�xy�+�|���?��f��Ĥ���/Q4�i�=z|�7��*/���.���ug��Z6��CЃUM�xݟ��oA_R�u������M�� 2�mW�z�,
��k��5�1��?�����J�n���ڂ�W{�k�ž��}/�n�']Ԣ9���۵�l�p�*����#C!_�qoiw���TpB0�)�ٹѫ$�s>�#7e�}�ڷ�f���$��������W8l70��e)�ß~|��1��N�����$G�ܽ���+Tk!3�!~����'{��"n�,!�W���h�<���ސ,��M�@o���0���:�j��&7! �$R�ke�ͽ�@���!�H��r�ݿ���h�-_��-�j�)pվ�*F֊p�F�`u�v�$?��m[��~ٜE�RB;N�D#�F�@�;���i[�Jӽ��5��oG��ĞykV�L�����|A|�}�7��fb<�o��vG
Gڨ}E�0uY��C�88��jCHO3���ſg�a���}[�����n����۲�SɎ16g[���$˅�;c�y��0��Y��X�GDkA�\Y4�Z�Y����B�W;���*��Q'*�F�w��=�ϔͯ�5�O�p�4lF%�b�e~���T�H����8c�䎲R��܉����^3�����^vk>������;;�x����+iOa�f.|t�H����S��ytˇn��E	�����M����Ux>H|(�O�P&w�0xW7��Aȯ%���akm%��:��ʻ�0��7���5ot��(ܥ�����R��Z�/5�̄�^��A{R�F���d���t�$h�i������ݜ���p��k�56�n����~��Z:ߋr�%�S�m��ClO�w����N()h�#7p�V�4Dk���/�Q��C� )��_��ـ�����b�\�E���l 鏙dDA�E��J�<�*�5���C��;
�"��2��¢Oq�K�{��3{�X�y�.P���������~L��*�E%��Pi�o?����h8��u)~�b6z����,M��]�Ÿy��흙�H�7 vEV��6��uE9��y�.��=�9"A+�}R�<P���ď�sSqy�����X*=K�������ɺmP�:���o��s���s��0_RIf������^�d'�}I�8M��Ne9L�T�k-"�;Aɲ:��d��W�|8j`P�S%Σ�	�qK����/��bv�A��
�J➣�d򑿍�)��*fU E�&��Jn,:��-Ol����=
��mgx5���ě�4iȲ�JC��?6�wΚ�c��k+�D_�g�t�����n�&�-o
ͻ+�����w�2d�0�aà�c�Oܮ���F�U�o_���?C�����:�Ӝ[�;)P!�W`���u���� �I�`u4_�ڰ�t�l�ȯ��6��<�R� B3�h����!����U� �x�?1��qȭ;:�Tн�IV��Ԝ����['�����tU��?���becs�0_���{��Wf8��'o�LB�7W���?T�)�is��'��v����xB��شxu�-��]��S��Β�W�`�b{w��	��Wx���^p�4�4��$��2b�ܱt�l7S%� ��+B���N٥���ȡc/�A)�Ydc�,��"����q�ç"���&��X��M��̚��a�m�;IWK�ixO��&-��8�ϊ�DD���P���m:`�3��ғ�t��@[7\4�a���B��O"=N="�D��Em��r���F�m�ڱ���+�R�t���4�ԓ
�@�N�ܮ'�=y�������?D���hv����w���*^��l��BQ��ְ����s��F��%�x�eX�R�lڇB5L���g��n�jF2���:�2LFKyJ����7m1n��
w�k�D�8�DȾ�5|�z屹����?#���]8��(�#U�9/���K�R��bY(n�����Ter�9Q&Xn����pk�lk����bHd�C�}8��c�mrvk�l�0dL�&���ʗ�:��i��?�{m2�G�F/F���z?��gƱ��-l��ݥ����~{?��7U��D��W��꼮6���)�$��&�)�����Vq�.����3.�K�k�̩%$R����J���x ?Ie��\������~l��$%�&�R'��l�9[�L�6&�� ҃�Q��{bl��X��X&�i���#k2��e";2	xzl�8����֩j4U�@��(Z�����4tnA�M���[u,�ŋ}���9�^G$Jː�kϪ����{�� �:�6�����qvś���7!�c��{���[!�G��}�	�O�������n�_TA?� ��w���?�?%%�ރN��M��2��	t�i���	����f�vX�����W0x#y�O�u:T3�ۙP�
U��\_����l$���#���x���i��ka��iQ�p�&������O�'v��I�Wn��"5�|ӿ���tȫ���M����o��U@?��jݷJו��[]�H�P�U$`.�m�lB�#��f�be2�}���z^ ;������&��\*�][�ъ�ֽ�zi��Oֺ+27�N��C���A�W����c��Zbd"�ȭ����n~"S��[R̽o�!8�b�\�� �	��j��P�~E9v��54)�ciy�a�*+���+N�k�˓sߝ+>��K�����l��t^K�h\{7���/-Yl�G��0Q�����D&zj�.I&�|Ȍ��&_s��ݞ��4 ޴��
_h��,�����}V(r�ڔ[�>`��蔆���A>zk���0n�_(�ْ�m�Q�q{���Eof��g�t�Ը����oe̓�>��UAC^�27�҂Ŧ�oȰ�h�|�{f[�H�=yx�j[[TkY�=�-�X˗�IR��ѫ�Y�[T]#<�"��>��H������W�� ���\{j���kΈ-��c1 �SX����+\��FE̜�ǻ�~=���t
L/�w�gaW�v�Ce4��A�S����W�������3=e���ˇ����y���Q�8�W��/��P���'��c Q�lQ�o�D���ψ`x��_�!�@jWC�W�y���Aщ�g�<#Ҹ�t"VW7Z�	�΁��蠖�����2Z���H��H�Cw��Mo��f�n^R]A����v�����.��F@��fU�~ٚ�,��V���`��������rV�ԑ  �{�'��i�\���W�!-<���0�O��v*�����g1�kIɆ ��� 4UȖ��u�~�5fL��y��i�2��p��{J��פ���������hH��0�2c��[el]�b�x.Ư_N~>-pP��ƕ����[N�Y���"��-�*�VC�O:b�^'E6�7���9�J��*�z������`;��5v�Mgj�����lk�2<-%����i�Or�������Wg�M�r�����"�B����H���i �Nh�����!V���	㴆8̐���⌤�־�G59�JK�3���;�4�2jc���YÐr��2���R��n�����R%���E�Ǒ9�X���aYd��b�?�`A��^��0[�ǈ�a�6.I���eGѫ�M���5��W"�&�Y7�ήl��K��A�]���E2��2d�Y����3ZI#oPE�F`���#x�%�Խ!���E��4�V/�Tfބ�G�a��٥���m�p�S�h)�Im#Cz�2�C�*�"�M}A!����;�Q��o�8��޶0�(��+��>�l�Oئ4h��ʻ�� [)i\[:'���m�l�u�xQ�����#bqBS&qq�پ�W�u}��
/_\A.��_մ!M�bn|��f�����u���~���ĲT�I�������7��Q�}�v)3*K�&�5�ކ|��;���X)��k�-����3���m0�d,�uW٫0�)���!��hF���c͋����v"�>��P�v�GN��dq�6� �5xCr�7T�,k�HD�b����3������I�^k�����DztA��.���C��^>��V����:�(&�f��o��q��{��A���g�a�/M9K���|�"Y�#"���`�� �����Ozy�GZ�޿=!�����)|�X�1��2<
�_۪�EV�<s�������i#�� R����t�|��0o���s�0#�=�b
�{��E�s��6f�aa�9��l�-���:U�1��,jZ�à��������뚍7d1?������^f�'��_�G�C�_}�.{�Н�_M#I�8����]q�ՓYI8�r	(�č#Bn�*Eq�s�Zhn&���њE��-��t˕�D���e���vv�Nyh�?U������Sd���[;cΉν�zI�>~;I��M֛f����V?�'��Ui��7=�&��V��3d�N���]W�?��� Fǎ����Ѱ��Owc
���0�_j�?]%��b��2�ц��(-+�Mb���m���m������zH��ӓ�X6t�~rA���*���5�����LLĥ�_��}E#S���Q�l���`��8bS�H;`�j�[A<e�ZsP��8�W� <M�s�-�^�r�7;?�k,�A�pp����.F��R&��H[Ӭ�vk:n�Ʉ�}1��G�v=D�*�]��)G�Kn���(&>7��o�2A����'����CpXn~V�q{Wf#HX	ޡ����K.6+	�P�X��Jeބ�K�a.PZ�$�܂/ki��AIa��&�ݣ�!��4�[\M���%�;'�����3��4���C�dpw���·�����]u�=��W��Æ�#��A�>sq~�5��o�+��j�xkL�cA�a词�4��A�Y����:�3l(2E��@���{"J�#Ah�i�:0�S?��H���� L!Y��:�F�U|��pG���Va�eJQ�'7��7�������7Z��S�e)�_Ң����f��Y/,�Dѻ�I�V�=~�%TɸV	�������3����R���C�[��"$�ٌ6�v�X�@��ݟ�ek�##�gZ��.���q�5������ ���*���_�)�>Yǐ��C�.�#m��n��!"�9���ə�fA�������e�#�Kz�K��N S�0�XD�U�#���Q߆�UT>}�m��*��t��q3ej��K^d��IM>��Z�b�z|�h{��:"칡�u?�p�x�G&���}�k�G�{�v�!eE`
dJLȎ1�g�RT̀Z�,��)3�3*h�Ei��u=�=�M�~o�;̮�V̇�X��-�P=n�"j�d���n�G�i*�σ��;W
eeU�������Tg��K���YF#~����Cb�ŷ�@�!�FC��o��d�?\'M��ۉ�;N�!r�&!���&�<Z�v���B}�#
�9��@�H��\��ձ@�S��WRD���<���]�����K쓾�X��KԌ���3��k��n:���S1��O?�����s���3����F���5&QU�=���l�O�(Ȏe,Fm�ҡT�c����^�c��i(��6P��`<�P:�����( cĴ4�*�ʓ�灨X\��̑�{�Ҳ�'W��$&����:Fk������D"���Tۼ�w�Hr��Y���Sf����
d����}sbB+HT���*8ʩ����{�Z���U� ���wŗ���I]�p]��+������d�4������XQd~��:@�K˩m��?�8�%j3����þ���uB�V����g�}���37m��'�4{hD��/���ξ��'%GF]�������O����G�hH�v[���G������ea�b���tCR���:�N���)��_�L@S�H��y��Ǐ+>�P޻�(_0������w�u����娴���q�1��Y��@�3�²�A�V�C�7/�X=��c?���D�.T~wF�$K�Z�w#���x��t=���`�G�h�k�#�i������ 6w:\N����w�)!X�^��
p�	�M���I��eڎ��{��p9IMg���֬A��@c���k�=[h|޾^�4��8�Y�#q�9.��
�%��!�1�V��������M���b�ߛ
n����U�Uydw�u�� ��ʷ��t���;ΉJ�m"�M6��i�G�����FW>�w~�c����ϰ얊���<���is�h�P�Ǥ��9�ٽ�����E�� L�4.�en
�ԧ�7�������
d��>)p\x�k�6�B�=u-�Y:�-�Ur���yW���̬>oϥ�BV���*DE��zy��B�
�Di]��U �`���%o�Fg�L���kL)%Li�����������2�����>E��A�bT&�Z��KA��%�Bwd�r_e<%j$ƀ+����ί�h>�=ّH?g�o���Yˍ�_��[����x�!���e��R?��h�E{9��.�P��jY̥��.��-���n�r�I栊R���Pk(9F�w|��-@h��Gb����|8�{=��Ю#�b���ڼc�#%]��))�� ��Qp,�K��m^<au������[�C�_G�����jr��zm5�����l������X�f�ey�>F�GRMj$�n|�q�H�B�m^����S����ju^��`$2j�[U��Y�~���v�����zB$�"|$+���� "�{���FCA���#��l�����,܎��X�l�6%�y�7��3\lܩ�~�)���G+�-�x�;���g^
�A�-�h!�F��[��0'��/��覽��,���Q/�T�w����ug��<X�󎼲Fe����]Mtd"AE��>8l���[��-�+)�h�]S[r� &T\��u�,��L�Iw'�ʲ���#f����O�P5ٮ�2G���3���C�,2��j���J�����n c^4�o�ї��d��e� �|KIֽp}e�gX�K�L�״N<D�
;�h0�zc��l�H��2��QpԾ�0��|g��}oN-��+\���}?�qQ������(cBBU�?6���n��8m>y�}��&�������C%�.o�Za�Q,��o\��-�e��Ә*���t.��͡RJ6���DEjL�KS��+���5s��.V�'��P��_���|[���<>�F�?��.�	������[��g��t�%�z�>vK#�8��}>l+�2>�	J��S�kP���F�G�kˍى�\؄�	m�;&{l1���o���^M
78_6g�Z���z~ �;����֥����f���kF�O�FZ	G�!H�m�@&�)����cN��Z"�4�^��05�q�����2b�����翲/�`����޸/P���ǻ?b��̚��:6/����N���^Q9�S�Ch_�<v��ID�t����w�x��JK��)N+�9 Yr���B��o;!DHb	�����r�=F̂c�,ʆ�T��7�%^HpphM<�����Cm@D��8���.�?4�q��ff/�m��ib��Sc�'ڒ|�
��Qew���xj /o[�/�A�>����S��m��R��.�xx�a�#Z!Nn�!�N�58���6�lU%����C0��-���X���%I84.�LY�v\ޞnѩ�;X� ��.��h�
���u�B�ڦ�;���<b7RM:���Ȭ�+o���t�`Yr�U��3y=�{�������S�!v6�N<��_X�����j��,l2D����X�5#�Ȭrz�w}#x@�;'�k���#�7�/>������G�����\3�n�fy���b��.�i)� ߐ[� O��/��ꚗy����e5�uU��Y�Z�Z�.��U)�@4e�eA���LT���!�[���<��v�	f���B֨�`R���F�;�D+b��f�nD������Ğl>oV�������L�&�/�����v��86׭&AL�b� �asdb�L,uɲ�4�z��8*GH/���f.���n�T>��DN:��$���uV�V��W�$K@�� ��<d^G׈6��3�x&(�X:a9��ܒ�t�������Z����*Pޝ������n�;u!x��9~�d/s]���O���E�5�c[�{��A엔O��h��V���ׄ[�l�Qܕ�id
ޥ/l�H���2~��f�H�<g�b�< -
�!h�rO(0.�+cP�(\�ź�w�i���[�����6/J{H{�dk�4�j�܋ۯ�<j���X�<��������k�D��%
�1s�p�L:��YN-!7s�+�o�hiÁ�J+ ��<d�)����ްI6�q�Η	�����?�lg�d��Z�Y�7�E~̝n�߸��kXm}e1�i��K�'�m��|�n�N0���ݮ��\O�帖�Hn�~��\�A_�&�+��N�����!h\��%���Gg�T�l��jx�7=�e��a���@�jdI��j�pD+��Q(�%	E��#u춣 �
�H�H�Cn&����TM8�H���c��-?@�e�{mٍ=��p»Z�Ɣe�B�Mb}!�����c-�>��%؞	:y.�l�u�U��}�a�Z;H��c:�&/�*��;�S�/!���`�NAifb�,,6]�"hq/p���� �L�A��Xÿd���}ƕ,A�%n7C�*$������I�<���͡eTޭ�Z!�t#���y:�ƞ�y���FZ8;~�q�h#�:�\�FE����<���:5Z%�RIO��܁%�sWK��.��]]ś\��Y���\k���z�:,�U#�N{��!E5	�.14� a���p�Yi���|I��lx�m��6�� R�����]�`'3+��侷�����y�����UN�`[)K�Arnl��,I6��d�mq����KN�☠�����y�3>m϶N�;J�7�	b1��pv�|K#t/��4|�`��#���}RG�94j�boO��LM]@`�Hrw�{��%?�����J����!��K��uJ���[���*iL�7�3�/�F�8�-Y�_sP��Y���KӴb�3a���=�<;��Q&r����䩳�5d�&�����#j��c��8	�72��˭�=��]^?�ݎGԳ�;%ѽ��bh���8u��E��!��}Ys
�8_�3ٓ���h��#F��N�+���"�'�6���h�K��k3����(�8��T�)&�y7J
�Ilx�ԶR�5Gu1��e���~ɭ��$
}�÷(�)2f�`Y�٫E��#4�}C�u�K�KD�Ma�O���ְ,�<�K�:Y�l�m�$�6"��0#�N�"�'I@�j���U26hZ��'�}CSt�1�1�nR�;��3��/����J��/ى|�[�?q�$Կ�2�U����i�J�3D����r��r޻̶�>i$�0%����j;6�$���I���K�����ތ��G>~�;�o� ���M�
��qw��m껼�L�X}g�e�p����6(Z��U��BGS(�,��8��R{�L{Y�?�|9�ҧY7��U�X�4ɠ�$�f���p&���o��!g��Lͼ�_7I�b`<7�C��~�N;��t^�7�4I(���\�T��\!�4���G&�K�&�#,k	v\��s����FNm��8QƧp/��+�A� �1���ƹ�~wa�v�2"���`���6z��c�6<�*O� �[��p��i���Za��.��Гߘ������� 	a-����]-�gh�7�]V�7Q���/��u����ysO8�\��-���n�$oeBe%�B5ͤ�zXLe־�s�M2�	�x8�^������v�{l&v�X9Rs��L���r�f#�Uv��ʸ����ߚ׭��h�3���u���<{\ᘩ�	W>����]��X\�
A<�-�Xam���*9a�*�C_o@#��6Ω-����(��I��	�a�9�����w�����=-`竨'݋;fS��oak}/�'{@>�'|u/����ɑ:���9,X���5�^rrp���K�~��%�#���-���7�E��7{Z�uH�Uj�=����f��X�05=����]}�>�P�{�D�7K��E�pQIW�F�Ϋ�zh�d�'���Ϯ|��&�����v�$/$2�f��ܼՁטq:L�9o�]�c(�1�E�gI��J�e�DB��#����\���)c��2���I2^��Y�-�=���O����g���ҞK�U&��箄�������bBO���^}��y5�M��eQ+4V�IO���^�/>oKc���%N[ˣ>�|�\���.�im�-�sNݬhy������`�K"-A���Z�2����_~^�E�w˽  "UbTb���c�E�]��z�S����H�A=��LSO��{�,˥;�#\Lk�D�z��=EE���"��x���6J�[�=���Pό�X ]n�3)�'���74�q����&RXp����=�G��AFK;�k;�8G#��w�^O�Y�-!�i;�G�4Y���⤉[�?w }i��T%Y7�]�RY�	yǾ�M��X:R6>��e�Ug���W���m��Ze�!mԙ�&@�o��*;�JC_����x��ն(�wƲ~d�I!�� 4�[SO�J؂�8}F)�}
(f vq����|Wi�����e�umEbИ���\z�iȸ�9�m4�V3�0���R32�^E��הK�����5�p'}��A#�
�R�zD��Ŵ�b`X����
��)Qi�#���q˅F9(:��<�ERLXQ9c{=%���@�#���S��!��g���>~�+%�mB�.1%=�������M�X6�"X?��4ظ}�Y8H#���g��Vr��u��ॅ��H��8iS�Z!�`}K|��������)Kww���!Ο��)bu��93�	��^�=28��f����
g�,�7� oI���ة��8%;���R:������� ���g��G�7?�^�L�,gG�֏\��T�հv�=uN"ZB�������".�*O>'�c�9�8�z��g�jN� 3	ALdZ�om�K���zNr�Z�i�Y��|�w+��T�����&�+��V�(�OJ3���am��1���)K�o�Z����[}Zz�z�������gw���@m�_�
%�K[+��q�s�� ��:��|K�$�'�9Wx�4�������Ӊ[ܴɠsU��T��v���516"SƯ��(�C��B�x���t�R�T��o��cB�N�۠���)�7�J4���h�K��&����J�TvR�(<��v�5�᭢e9N��%�tX���e�G�}�����u���?�c>�������sn��
��1�^��6_ށ�ǈ�@�%�l(�c�p�bk�7��/emx���[M �=�����#���ȲcZ����.��İ��3�v���W��r0k��C�J�����n�:��_�"�>>���+Ү1P���P�{���
�^�5���ܘ�����e��*��}X�N��<����{����+�y��h�x���+K�O]t�.���E��w��[	:9\n�����)a�����[�#4/���j�kh�c��b�1+�s/�6Ú���߭,3�~��χ����9
;��F���)��Q�u �A?Ty���T�c��w˭��b��D��vX�3�|X!�[2�t��'����d�@�3��%�QD�uM��V�e�h�7π���j	�1�Êm��_ � ?����F3R�O����3W@�Ep9��Ca%w�{�p8a_5	�Ѝ�e
?�v�W�,!Y(���_�'V�Qd2\${�d.K�q~��yQ4/�]���Zs�4���[���3t�}�Lu
Y.�m|�_<Ny�p�&���9���s�Ȟ�;H?S���HB��_��l��� ujz�ƾeT�6^��ܷ�	橿wdg���^9����6�M�f"�EիJ�q'��}vaY��P���X��)�M���Q�["ݡ��e�F{}����F"���ȴ���:		�(�cZz=I)�d t��X��?�ʼQL��D?�ylQ�fQ�{\G�)��c~�:: �	�K��V;�ȏ���\	����ѧ~>��E��5ߋ2�>��𢲻�p��V��:������3�~�����f��#L1h�&��Ȭ�����?Xh�5�xt�]%0�tIP9�մy��o[�mV!j��ȟ�U)�M�g�f T����X:�����-F+�G�m�ͧK[��6B�~D����x�|����;��0N��t���湱��Ǝ��=(NVnz܆�����y;�����a	�|>�1̸���,�)u���TU0���ɏ���N�����]О2�su��-�G����v}X�{�Kޢ��w7'��p��]>l��\��C�4��p�z�V��h!�.Y�ǝȣ����[쏅��cXK�7�P���H�}]fA���d>M�'�΃��֤C��8l��&�Ӫ[%��>#zx��u��8���h� .~��8|���1:=)�+�����9}�C��]�v�JW÷�KY0l���>��A�AX\�����{�d���}���Q�r���?���T*����(��A���K]��*Zr�yW���/xza�S��H���VM�o�����U�Z՜%�8�9O2�Q�����U!xy�D$����suNk\6��IJs�����Q��lK�G�b"�_���B��YiU �=��S�䮼��=Zʻ�"a���oA� )B]�a�.�
_u���_ڊ
����X���ۺg���{c=H?M�/a
ML����G����p��݇U�R$4�3�,S5�*B���'��)����
�/�pd|j�4�A�#8�.|X�2��O�Ʊ�K�NK�_�_s�o������&"���U+�.��|�Ge5v��w���w@��7�K+=�$��̕���
Gp�	!`�E���ǥ5م8��fD,-8,G��DC@m��D�/L?�Lع+T�#��U�1���d���6������{k'�~&"�6�=vC��ٹL��"vq�9۟rׄ��&�|�),h�e�2L�6LW��gU�dǶ%�4J5�2Q��(:N�c)�f�W���|���'�O�&ߦ]bJ�=1&�Pۤ�h�����g��h݆k&�G�/vb�ڜvEi���(o���)�9;ݻ��AM��OE�E�.|�%u��� �ҥ852��ж×bh�����A�����%*7�T}�K��]4��?+��X��}���D���Z�B����c�g���M�R�s����	w�pr����ݴhֹ�?��j�]��o����w� ��L�o��蘑e���/9L�5��V� ݝP2���F�	X���M�����<p�Α��V��d�6KJ&��*�ڲ�`��eqW( n3k�q��,�}�{�O�L}H����ׇ�<~�R��1,+�R�;&f���h^��ߚ�m�M��ڎ]�p`����j�oo���z ߹�G���F�:li1)�v}��/���8����	K�B�������bɘ9���{��6Po�I�jh^��إ(O��g���`}���J�T�b-m�xS/�p*:J�s���_񫦂jqZq㊻���QzKv� ����t����+�kO�"�D����^@������e1%���s���ݶ.C��>�0V�o��?�8rȢVC��Ա���94�6�n�n�[�y�,�S��A/B�����֨2[�Ɓ�$#P�����,K��V_FB�B� G�G�j5K[9��\	X�X���Ŗ�^�P���p����
J�*9�榿�\s-
n����r7� �͠�����t��!�÷l�}u{��"��G��*�F2X}�}��s�g�E��_�"ujh�W�V4f��<Wg䥶���.������a�Ŷ�ñ(��]�0o�1<]�n��b�ɛ4�7���+ �T{4Dh�3�m��h>���;��Sc�H��~�`��%#-��Z����������Z$b������ͮ�L�$�/� <�^<�[ۙ ��/V�W�Zvw�w/��׵T����a:�2�G�P�1}��V���yb���~��?�t��[.yO���g�y=�"��4��Pަi�S=%��(���V/�~�%��/Cv*��#p�6��p�k�����M��޼�㤫#�,��\��	bozx��`�ո��o"�C�I�ߛ��TM����5��j?�D"z����z�ơHN� 6ҕM�Ɣ=Q���~ra	3�֦�N����W&���6Y���̓\����[���4�Dߗ �!*s�a)�s�cD�d�s���ո�� �@�5*ʃ>�{ƕ�B�ڥT��q�oѵd6pf�*���s��N_Ew��eB�f��~YԨ�B���}uu@x�`��zq�A�U�����I��,��������&�|�V��5Ą�e���F�����G������ի��Qgt����[2�C�m���ݖ%��
���a�M�6_��d)�'Ä3焵��O����[�od��-�\R�(S�}�����kS2���	�p�8:�[w�[��\I�c��r�I��>�e��eT4�g(�]*��݁�A�*���7~�&��M]"=1��"m�ط��5�V2Pa{O�6��V`W�q2xӀYI���i=�L��eג��sژϷ�qj`ͯ�a�3���æӜ�FW4]�E�+��,@�b0Z��"��knԈEՕU(o���m�_&�K��M�ki�����X�[�6e��ӕ�]�{�|9,Ȣ�s��gw�b�O#s�Η!��+�6�V��4������]�$\����DIX�~�o�:(D�:�e���J��Z��q�i�|:�a�>�!�fK�4���*�<���0�-L@P 5�ҝw;R~z�U���e����`��[l�)8.�$� �r����ԋ����<��^�e�n�u���O٤b�&�oɣ�d	K>C钙a�r��F��}F����Jm�����^A�� �yCk�
��U*h^v�G��_3#��)%⧌@lT$l�ߍ�t �&d�ک�G�:`i��A��c�o8_�;i��OQfq����Dl�g�L�Y������#�\��m����5d�t��]ǮSm��|:&�'?��U|�$��3��L�^���환�B�K�b�	�8�g0�N\���Z�t�S�BB�h���̞��1�M���p{�Q�	�"��s���Y��Cz;Q��2|��EP�gB��FW�a�&B	�Ȁ�bd�ˁyS�<�pvp�K�h5�ź������,�����cr�?�G��%_���Vo���+�380����A:Ș�V��;��*�\�E���s`��[6��}|��T��&b���`��A Bx5������c�E�o�m4�i���$��⑚����%��ᐠ���l����������'R���Дs����b� �I���f!.У��"�%����SBi���A���Y[5�Yv��O����u{R��q�߹P�&]�$�W�?%�?W�%�m�*�B����c'%q��tMqw��?���$����K��B��< �1p���J�1��xb�-5�ĤͰN& ������G�k�.q���ye�a:%�Ʋk���$�mMe��u���Ũ{�|(�����xŬ�]�b(Ŧ]�Y�	F�	7��#�P��Ԭ*��l�vSS����s'?�&��>��Bs���1����r�;�X��{�b�>�J�pr��r%g/~�ڬeE����>5�mb��T;��Z�E�}��CC8�ٴK�/!�����9$	�J�x��bg�5lo�>Ծ?b����~�͖5��+��Q[��Vi���q�:h�ȉ%}�T���kk�Bo�_o	�ΰ|�4��8A�_ �W�����{�?Q���܌Q���A���N�C)b�$�ո��p�_Q��ƞ��[��x��ڳ?+nx���f|�q�_?��Z��v�rܥC����j*b����v���m�9f<��.�;0�xǨ_|~!N������+�ŏpN����X�k|�WJ?�h뭏U�O��|���d�|�%JF�k�3�n�/�ޤr�N�6��v�s y�-�
&`Ż�s\K�C�+ͺՃ̝�[�!��d{�zS�V�¿H��\}tF{�˘Y���Z�!U�_��{ʵ^�r|�ԏdNS���ٛM���߅�d��e��j�/�?%�D0I렽|�Y�t�%Tr���}��j��OE��be��Q��;��A�&s�@�z#�^0��Q�R;O�%�N!�l���ӒV�HM��HԿ�ژh��^�K<��.���+�[e�W;-�a:�d
`��0.:O�E���&~��]�U�,;���.|�.;xxe�-Y��/v7���M�9���q��Q�D`�,� W�ul�e� v���O��3Ƒ��|8���e�Җ7�:v��|n�t��SsPw}��|-��/_e��~��|�����sܜtg��4��M���6h���WB�?2x�}�Vu�Ӌ<�׽C���� _	�<�O_��[!�4���yK4 ڸ�z�:Z�e	�H0��~[XK�9ZS(�	�4�F�U�%K&jڴf��`&�ɷ�۔��$<S;s��4��Q� (��Ds�0�o�l?2Q��j�U����tK�5\������=\�m(�[��ه�\�����tB?Kyg�
F�~��~�s����"�kYT���U��՞Rs+�;5�6�*���F��!{i�� ��Y�S�N�����������E	�Xp�����-?���\!}b� ����DŪ�=׵W�����尤�����׮�G7�4ʖ7�!'���yE� ,�}��&�܅k�?��J����4:��܏�e /���U�<�12!T�	�6���*t;�#��].6k����Y���fw�M���b�z�f�[������6;W�,��t��ޜR�,7�&�!Ƈi1�Ȉ�O��|*�рio*1� ��U��W�w���+Y����C�W�x�g�T�:���[R>��SU=�Ъ�=zR�8��ɃhK�a,蔱�*Χ9�[;���c�ø�_`�l��Fn=�;��+D�M�]x���@�3���0-G� ��4�P܂�e̷��L�I�A�N[	!l��؛�!���"q�OB��a<A-�_�8���p��ˁ>e"�q�N�MX1ᔜwy��iq����	5��	�,�$_�2���1	eܑ����ex�����W����F!�Yw�5y���Te�L3�k�>E�����~���m\6�q"�х�`���㤓�.���U!]Y�ɫ����w�8lm-֝G�lDƃ�0;��f6��O�����3���T笽ETW~��
˞��C77v�1"� ߗ��A�"���S݃u$P�5��3b�����Q�g+��������@��Y�2�d��#�:S,-�HnA�
F!,޻��R+%�f�~�;ڣ���]��KK}�K��~�U!,�B���r,�Z��hr�7�V#�u��6he��F��[Ea�{�U�����`耜GِVٚ��hu�Ɗy"��H��-��}�X���%��+R?�wd2˩N�����s/���U���Xw�q�Rlh��4��k��a�E
�����ZE�MȜ쨸,�ܟ�b��׳6J�0���2�NAL�!���`t��!�)I����b�Vm%�} Q�'�-�n�Rp���][��Cl	ɳ�
��:>S7�����`�5t�I�G��{�n�(�uH�]��wPr�̡�bB%���\�Pm�"O2��OR)�i��,��"`Kk�&�4	S��K�X���n|�>c�����Di�T�ժ�Ż���	cXѮ���h�1'$�������\���m��^����?:�+�#j毡�qeQ��L+5<Q8 !��p�_�*5a_�E���x�������-3��p�f���j���aBxk��ëi̬�s ,+C��21co�������Yh_�������t���]�`�����f����/�3�z�ĩ<�%X�)��F ��قh�i���PՕ�S�P+ ����֮2/��W��M��P�>S[�iĝ̣��=F?6^zd�-�8Z�8T�W�vN:�"of\���phl�:�a���}91M���"?�73o]�mT��_��o�І��c�(����%s�32�����!`�7+�� �I�M���?��t��؊~��b꽔��Q�F�~�eTH�ж���S������)
��)�ojJ����[Dr��w��	�k�m��!�3A�Di�O��.��WDd���+�B��2�
Z�C	[l�eP�VORk�l=���6q�۸S�X'QMBL]������^��7#S����r~Y��!j\eq*vY,��GOoy�}�V�7��5v���E1p�� U���+�3�Ϳ@5�;L�}�z�'b��+���_{�`���>	D�ɞl\��+W���"���C+nT�_�>����Wr�4AAF�$�W4G�ej���{��(:�K�)��^>��}���j��о�1j?7����I��ۉ��E�� Gkן�H��X�m}/8(�5�0�B�߂�B��Ԫ�R#�>(-U��&�7���X���K��_4��-t<s�iB��\o�À�Z"�2�I�K�%���J��U�����ky ��=��Gҕ�ԝk=�|�ӛ���`����"���eJC�t�%X���\ӯ�Un�(��n�.u{�ઐ�wS.f���;@�9��~n:����UR���d��f�M0Z��^?�FX��j�x���d>c�Kw5��Y�tEk?~�j�g�+aǧF��ju��k�W��p �pL9�ŉ3�Ƃ�f�MW߻Fa�'��T�/χ\/����.6d��K����C���������'�p�=�'5u���sB�"*�Zx"t��l���$>�xzA�o�'A�s=�G/�;P���eɰC�B,%�0��8�+��LQԊ�98l��\�l���5+ ��i����e�+�	�7�x��IE�f�
6�!ċ弹Z���P�����M�78�=���h=g�����7�-��~���	bBm����iܱ�jE��>ׄ��i+cMf]WH�tG-e��W^1�fnze\ �?vp��iO����**��"(� ��@n�;hWV�Z�յRx�f��/,���7�aּ��ok�_��2�Q�+Z��jYŰ �h#F�(���0���C�`g"2��ސ���XV�ro��Y���M�,$���{Q�{N&�7���N������'e|�@CP9�T`����%��5�>j����Rw޹��5�c��Ts��Ί��͌'�_M�H �#�Vɠ4'�j�z����2N��S] �t`��I$,�؊AI����_�xVGw�������	N�;y�<�yU-�D�zy�#����=?`0 }�t���?����)2|J��:%1̪���V�Ӟ@�e��WC�������3W=y��	<�ɯ&�JϜS���S���ha^���_�D���ل����45���Di�Q����/2�}+6a�0�f����~��6l�H8#�wε9�+�T���~�y�h�s�a�ܰ9u��:�����rG	3JM�]ռ[,�D+r�}+v5_���>����q���3�Z:):+���~�K��\ȃ?��_�Q;O��'�:�F�]�J�#���m�7@x�"ET\a�P�,*�L�-}������]81�<V�����d��a0[6K���?���m�n�>}�0���N�I�-�I��Mo~�O��S�l�2~O�Mtt��|aH���d���n��������>��O_�d��Jm	s6.�����M�z3��5�d1����1E=?_�V=Z�g��4�e/��1�� &����Z�U��Dz>����@�����|�3MӬug�OƬ_��� `����h�PB�s+.�Q�R;��?`4_�@�')	����S[ȵ��ja$ G���5����YH�	r`�۩��#���ŗ<$��#b�{���B|e@��i��u�U]�j�R�C����}ejp@��j��i�p?t�q'FXF�~��y��8(C���v�{���b��7�z��ۄ/EB\��.��[�c�򀜫%Yy��	��ԝ�x�2�)%�S^�@��̎QN��a�e��r�aݭ^J�͇���<�s��^=�t���A3�'#m��4:xg�u��q�.}��d|TY+�r�Q�6Ƅ{.5lg�I��
���_q��m]��]ؕ1���¶&�(�zm�%n�h��ؗ>r��p��l5�6�Z�B��k�	����2]�#�ݨ�*����*�����ŉ	�'ԢY�������8���z�R7�Z����iJ�	�Ma[y�g�����ך�����e�ԢvŨ������dsZ飝~��Ί�*�e(��o{�.��6f6N���[�!A�z��Z��M��1?dm��S�6�O�~��Qt��ZO�R.GBU9<�c	�nC�m�*�睟�~ӳ�/�=l�um5|�}��<E`�n^�T��a�y*0cUg ��죲��r+͸�,��Hɖ�l� �������P�=;�l���Mxo�Yٓ��egN3����O��>�g���ء��ﺰݳQ�OK��$y��(CE�nmR=#]2#^��[!݂�o��<����JȈ�LzV��5�c��s�� z�k��m�x~=/��x�-8��e�4��v�a��k>���|�a��*�"�����J*�O ��(�R/@\������������!����D1d�O+%���䶯ψt)ٖY��I�u�vvڔ��q�mW~�lLA����P�\�
�O���i�p�X��t���P����yD���i$]�g͔7�2;H��y8r�S�v��@	M���G?��Y�Z����8̗m�4������Q�Q�����"�v9���F�M^�;c����
 �	�qZ�'rr߰Y�9����M#Ja�~+}��Fm��ܿ�m[z>�zi�*���&;>HS�e��L�U`)L�k����L�ߚ:��3]7c�G�[�q%���ʨ^F��<s�8}8g,/;�� A;�z�X�'����#[4��B�C����'����aT�=:��k�#j�a��׭�����7�_KtuX�Ϡ���T7���W�q�� ����-V,����(	�*�F��t���w�f�� 8_Z� 7��4�-�x�ַ��}��f{�1���+�0n��f�q�^��)��B]���J#���A/�v��O�Ӊ�n;�	�IYkO��&<�f�q�I�p��y���s��T8T����%]����;�����UD�>�%����$���n�C�SP�NA��A�;�k���~o��?�r�yf��9����h8�`���U�Fg:��U�)'�_?���B��E��$�����nQ�Č�V��Et:�fa��{j��k�2���u��S@v~|�9���vZz��9<s̪I�������u%󃥐��CʩԎ�=&�@�[󠊂7�O}�� ��
�\z���hU�̝a�Tb1�)��}�4�Zl��$��Ky!��vq/,��Y>Hv�9�)ZπzX�C���B�M��u���c�@(�M�)���s-9m��q�V�H~׾�7��(��k`���Ic͇���`�T���kM�beP�@M�yH�V�&~.�����q(P0V��%*�1=';�y�p��%�d�U5�	�C?�W�3��6��7�.��؜�F��l�QR�T�Jag;Zӆ������|_SkǅS���JBV%�K����"WL{���������3%��|��.�v��,֤���Rg��S��	�yVc��P��Ƨ�WRe%O���Ԫ�7B��Q������5Y�����2ʞ�^a]�n_)%a����ɤv��I��5����m��j�YwS�@���n#�l���Â���`�6Jq�~cѨ��ȝo����,J��a`��'[[ķs����)���Fl�j2C�mתו���L���J<g&���g(�X���Ϯ��^�]۝�5��^`���$7���,f呔w�F��0KvE���X����ͦ� �ke4��n��'�{����ۄ���ӎ�-dᖸ5c�:��|�,���w���k����U��m?��V��K��(��zx��?A{vt�3�%}Ѥ�3W\�l�����M9���ٝFX䨗����2>�L}	���u�c���c���T�FO�����[+�&\ � ��>@{�"���y$�	���)Ž�����G9�1x�=.޵�9���	<�vo�U}��9/S�����i�!�yHYM糾Ox5�A
A��E����x#�oM�Eb���uL�wj���笠4^?�Q���eT|�A�G���:�ޫҒH.��~4̏k?%m���u�U:�u`���H뫣3��ͯ�Z�Oo?�>_T�y?#taT�e�D��od79@�AU�v���\}�EK%�n&ڎ��K�2��;vm��g���A�n�#���A4^\Dhx�R��Ւ���g��Km��Q�΄�^��y�x���V����$j�\��.�ћ��G��2_4UVd�54w+>��W�Nv�_����<6��������7d�ٝ ����b5���\J��z��Po�9F.���V�P"s���x|㩟���Քg�ri��)�B�^O�g�_����#y��ۖoЕ)�h��}�J�)c�Db��b���t�hU/��OnfsC#�ZjZ��;��̦.��>/�U�D��8�F��U" j�3Y7m�1o^=J��ׯ�xs�L�D���"�!3|˷z�NjѺ?C�p���ZZ;�~�[��"r<���*|+#Nx˄�L�O��u����LPѢ���v|��?{2Df���2- m�G�\DQ��ok`ա�ʯ�Dc�Z|ь�^#�m>u|���Gb��q�_��|$ꩅ>XK{�I��㵣�$�/6�$ۖ��0�K=I��q3Z�g��2A��J����Sg�|�w��IT�A䈐� ��w�]����c��űO�?`�z`64��sVE)>Cʭb���a�ԟG�>�|�h���5�N�vLu�o��i�~yR��bDN^l^vmD��F}@�+�Z�x���I�@ԙ��� ���a�zb��Py|����Z�x@���[�wO����H8�e�^b]��b(��5"�R��]ux|{v�&?J�������^G���_Ӏ�F�q����vP�r|ٴ哀l	D��6��
0��b9��3ͱo�b��P��04^�h����P�����_i�"
��aH�:���~�)�4� �d�C�t8R��<�f�#�q@J�0�{�����
,��Uj�����Xph~
�^2��S��2�o)�ѩ�{2�!��D������>eYXğ�>�D�>,h�̂~A��V#dq�Mh�hK@B�w���v摒|:_��5CE��>�m;�M#�3K�U��AܞR@����B?�����+�(��
��笊��4V��G����DɄO�����OʯVˁ�LH������kZ�עmِ{q|V�<�R�%�%Ҷ@[�+�����M�H�(;���wGZN?�D�l��
�z��$�7czEyw:wl+�/�������m��#�_�g�a��9��]���@ꨌ?̭�"	q��
:j�h-C�DE��� u|�Z(,7|X����T��&�����������y�i6��ޖ�]��|WY�,�^�N�
�s)��`��xT�(�"��k��L��R`m�;M}٩����G%c+K���Tz����,��X������ǎ�i���]gMTYt�5��Q6�J�/�Z�t{ʰ��7��e�j����E�P��y�S-�ܧ�Ʀ�����Bi����
�׍6���V�m� �:�[H�d�1��6�D}ѐ��gA�O�ړ�Z�JF�?@��	�E&��4y�9R0�(��&�M#^fgX�5��!s
\�?�L�����ߍ1g)H���3�L��F����R�m�_LM��#\ O)�ڄ����mWVp+`�ߐvn�*UO��L��gD�X$!�õ�G�j��c�i��9]4O7i8�/��5M�]� &�Y����*��z�'��W�l^���I{�0�E�t���2%Ҷ{�b�f��G���r�
��\e�B�%~���Z�ax�Rg���&u`�|���%���~��x4H;�g���vB�C�UT�ج,�._#z>�*�m�/0=���QY��&#n�F5���`��}$t�s���7��F��e�b�TקB8(��Fg��@�(�)8�4-��
%;����ˌ�?7]H��@+���,���Cpwv�����m�В7.*�y��q�6��ؔ�藉�J�p��M�V�)x�n`�F�IZ'�]�?/�	�V1ԝC�� ݧ�F|�B���F����[A�l47�˽&���w�Sc�[��Smx���<��\�uJ��9���t�y�2����#�[wP)A����N��)���"���&.��#��iz���`�dv��%�'�ئ$��jC�cQ�f����l�m��(0�n�/7GS�K�d޵���0�F8EbP�����-�	��+?I�p7�@�fO����d�5K��ð`��v�D�cK��<fVN,a��=#Q�����seN*����R5���@��L�N���'	l̋��g�V�JU��i�/[A�_��H�K�-�3ּ�Vq�!�h���C޷&�y�W��*	]������72'YG�+y6Y���*��"�W6~��7k�b�z�M7�(�a|�uv]z#����Ǚ`��f&�����`Xⴧh���R��.���ň
�s�:�.� �:��%��m5����۔�qk�ʒ(�%n��;ҷ�\�F:]�������jϠ�=*��[��A,�J��8�Ð��[���Hc_S9h'<�_�)Eӂc�02�ŏdR{�vW�a7=���� �~��!�e=T�	5��7����3�¿�����#&�|��W~�G
�ZӢ�h3��@�C�vJ]]���E�{�����y�LFM>	��y�N0��m�/�Ħ������rX�c�~	s~5�{L|u�P|P�C���z��o�D���Z�����<��2+ZK�h�0Ȟ�*��� ����g"ъ��bh�����AbYX�R�qJ�,mt�`9�f;��y���N��%!X��.cXq� ��\��'q!Ѐ�x6H*y9���#��%l�^o?�E��3�:l.�l�[�ȿ��V�*�h|y�����������[>���!���^�Nsz<����X���WK�nB�,%(}b�%~�K�!�95��.�{� ���}��prG^�e`t�6�˯�{,�r��?��q��^��,�8�t�ޑ���e�_���9�)�n�*�K�%�����+��ᐮt�ֵ�_Y����L}���8)Ǚ��FZ""���6=�m�
RK�ݍ#�̷��B`gAknZ��Ú$$5�m��Lhn�}X��`�e5����O-8�NOV�����×d�嬪��R��M��K���^�D����;Q�+̐����{��U���?�Ǒ�F6����8~'��N����q��^io�|��XG��kۆ!P�uP���n}���辺F���{��/=Y�j��(��r!3��o��ד�����<�K�9b\6�-����t�y��@FPlg�Cm%�#��OI���w$����qPh�JN:'���W����`Pi��܍3�Dj�g���{[��R�W��>�eqFɗ$R��\�5���,�z��>^�}�xSj)���ۃ�U')=6�"���RNa����#�B���4�Ugf	���H[)V^����-��n���r`�ltٲ�m��Y0nOr2C�n9���n��em-0.��V��kѼ��[Z�.� ��c��1�a�Vb��7ڗ�������KI�ks�iN�M�D�PR-���Е��Ȓ�F'PQ����"���S`��x��ZA������e繦t��d3��_�i� DHe,�Nss.�����b\�$�5�Ϯ���M�x,����29�T����y��ړ�ש����j��	�x���vg5?��{�nk�lb�EKߑ�̩�+�����,3��ZZ}��%d�פ���0&��L3��|,��ɳ��_	�}C���Shx ��'�솃����j��E(]jM6+{ٔ\uP����[,�֟��? v�-�ל�`��d�M��HUƤ�p6l :0�ْG��#�!ZhiV[�C�O�+�>�{}���zK��n7����>6�?M�U.r�Uj�/䌴�����U�b���J�F��v�C���!%8�<o$�:�E�3�9�vD�d�!X^4�_��΁J|�w&.U��Im�iz!?�\:E�&4�L,R��ǱG�0P��6sQi`���oӉ]���hHn�:S\f���a��K�v��n�d�5q�_lC>�(Xx��@T%(�����`�e&�CR˺l�6��g|�LnU��+��3v�J� �1B�o��Yn�6o+��^��0����ൊ�^ ���0��s	X�rC��;h��N��ԛ��X�Ds�8��#�pb���.���9��]I�Ȓ�u:0S�)|��O�	,/����1�E�,f����1���_m����$��t�=!��V� (�j�}KEb�I�@�P�^f4�IhӔ���gd�������|6�� ���&uH:a�~H3)B��b�v�ͨc�z��&B:��b�NkS�e�_�J�C��\�����V��"�=�a}2�q������T`��<d14�e6C=�C&�E=dG�j����}���4���Y޴�)���KjD`���Ĩ�*�;�tc4�(���;\T���НLE��'�
n��s����s#�d3 �������8�S�9|�F��'��%'@TA��x=�����10�'���6!8XF��j46�ݖ@��)մ���S��h��n86��Y �U��R�����a�����T��!���M���㇞�1�+:�P��쭱v�͋xؿP����(�����Y�0c��2�R�=W��i2�7��͗��L��:�P� |<W�w��l�9�Ζ��-��}u�93J�ߨ���>ni�����E�k�nY*8M������\D�S*�ҏ�wtdNl�r��e�BU�^�^�.�_���	|��{��o���R+�L�n}��:�5��;'_JuF��?>�Dz!�C�_���݉ף�5Kե�Uz������"�w��z��٘g��9�c�Е�h��7|'I��vs�e�����E-��/������E�J{�C���=�I|qua��i-�^1��pk��Ȏ�[TM����8��6f�~ʤ½bk��R]����ap-<�����vr9sh�*��Nm�:>�-	]#�!ȶ�)����*e�ǂ�n����F����E��ԡݸ�,ˢ��>댑��lQ��lo/���ԃ����	Ϋ���;F�'��m�.�
��f�?9��n��ꕴ*v��Gh����ޅ	dG�	��7�����K<���5����\d�e�g�փ/ّi��R<�Q2�-3P��6��8J�v�ֱz�N�A�k|�'E1Ւ�d�`׭��C4̆�ۭ��1�@�bI��;�n���C�4�s΢�s4�9��M۝Գf`N��t����i�_�o�:.�����f�2xܾ��E@kjehj��������dkO��>oFM��o��6��a~x�0��!0�[�6��{�K�����g��bF�=�n�	�l�nT���S+G"/�za����g����h�ů�>���B��O�=���(�B���G<;�(���"�y���N|Г���Hg�����w1{DS$���t-�8�Q+={ن�)Կ�tW*�)����ݡ�E¸=����}��p���
m�p�´�p&��?8j�+o��/`�ԛ��U0�|ZY�M7D9U0&=���a������k���Z΁6π�W\;*�ԉI2<��O����{�q��K"e�	G���AJ����(�@<Nf�&���'���+���]]�� ��Aٲ����KTp��<;8t��4&NZy�r���b���vY��ƺ��!b�Kv!途z��m��X��6�XP3t�=��`��v����q�j��¼�%��Pn>e��N�G8]�.��w�@U��ҍ�/e$��m�U�ފ�6j+P�n�65��74�%����}_�Dh[�ͧ���&�����E%��J-��j!^�rS�9ԙ�G+�k��5�KZ_3�6�횴�8�χ�,MV覒b$Q�4�9�Z�Vk:��=����%E�Ɓ%g�Mϖ�;��A{�4�����VY�ں�on�l�/��p|z����7��ٯ�6BV_v�c�	�Mc��W�"y}ţq��{�9�[�`�k��%R\!�Bw�A���W(����j��z*|]09Ф`��f>��ՁF	���n����y�=���t�W1�њqB��b'JHJP<3{�H@��^�)X1,��WU�߄>�u&1L�?���;R��ɨ8� ���qH�C����j ���=�M�=�(�5���*ͥ `nS|3��9�5B��0�`z�<���ON�f���@�y.���E�X	�U$�����&{=U������A#M������P��Iͩ:��Wa�6n�(������ht����4:�G3��UX�F"Z w��}4�~y#v3�k�����2��L������#����ԁV�+:���]d���k�L3^츚6i�j+�۴9J������n�I�>�%�.(6�1,M$���"1_j0�AiO�J���ґ�`�[���d#VLC�ݶ�cZ%������w�ƭ�fA�eW�As������[�2B���c�]��Z�6Z�Ғ�hJ�p[$S �p�BF𩸉.t��O1���*����=���4"y;�C�!)IfE�[_U6�)f�����[��F]v�����-U8�mp�ƼS�������~`�l����*-鳹.r��s��,`��$g{��Cj�NU8�>H����7� m�`!�i�*2'o#M�C=Ιg����Ǆ�3�ϗ��:n1=�|����a �~�v�����,X!/\ҥ��� ��[q�娽.�0EW�;G[-i�+8�-�kxQ}sJy@/	$!��ZYџS��nY}�!�U��d�w�Rlఋc���n���G$Z���{uoƹ������2S�J�E�g������D�MU��#��B�""����I ��c]�H�Rw�>��K6�Hd��
IRHi�b���i��藈ic_�Z������!�|3m��@G�1�D��05K;|�SO1��Ͽ?JF0"�����Wӱ}��'�a6ݐ`�T'��AiRnX)����B�L�B\�J�6���8�Rc�x�ˣ���+J��1'�̶t�(9�����<�}W:�t�,�Gbv��Ri�	V�x̵���`��E$����=Cd|	dS����B�w.�i�3����Ki"Eψ
5�¤R��<&����5��N1�����f���K�m[z����ry	�Y�ZsIdS��PxM��i^��|��]h1v��K��,v�א|t]	�3��|2��\2��DG1W�������_[��z��BB|j��3��]�� D1L�|Ɇf�q�W�h��a��E��2���D��ӈ$�6,��>C� ���a�|<�Bt�����4	&���Z'��.�zG;���V�pǶ��>��`M�������� ��1�9�����Ӈ��A�`��Y.+��х�t�2sb��Kn-(�w�|-N�����s-0�*R!�'f�"<�G#��D�-�]�&��	�!�$�a����k�j H�Cݵ��qY}�ƈp�w{����xI��ψ�>�یt��+8WTZ���^����H��]�����$����Za��GWWPȤ�2�����%=27{Qy�%�"�`�T�s�N�ϭ��٢k3�����I\KvG>��eպ�d�Q�^��D/�$��^�o�궋��*�^��wա���>[NC���e�����=�l.�K]5��T66�ݦ��e��ҽ~=D��&�M��Sb�����oę��y(�G>�*��<u��ӣƅ�E�Sˍ L�4�����Kh�o�������I$B1��וj\�>��Ǎ�!y�~X�6�m��~�xA^vZ��?`)�7�UY�H�-�:J�hg	뗄�"L�h�<8M-��P��;oٮ3)3�J���[��݀x,&����h���"tک��N���'�7a�;�p>�I6�x��Ƀ�VJ[5L�M���٢V.���}�\�cX����
$���}
@�=��am�/	���©Ce��%�J���F;�ǳČ�v���ܛJtř���Ȭ-!<y�|_-D�~���xA�4��h�n�:o�"�A+U�2_��>������忁�t������X��(gq�@�=n!���D�^�N��fIK����D�2�'sw�Y�t�U��5L�?x2�z�ɝ� 3\���[�����i#���=���0h���q��ߥ����O`B4H�8��_Y�������\݅NV��M��ػ:�A��R�`!92��ݠ���Mp�i�k���m��x-X^^~�g�;�'�;5��"i��9c�.�3���/��A?2�֙�ԒڄDS@����mQ�m�/�9t�J^Se��-|�?��_Ǉ*�{���0�v� Qtl8�.�ܡӼ�jF�5��5{�ܝ&f[֝�ҙm��K� ��~�h>�k9�	�XImo�s��w�^��5H���t���k^����D�6�wJ��� ���0F�mqX����!�\�8?;|D�����kL�y�d3�UYs[�YVy��v��5��W�F�4A;b����\W�ak���^H�pj :�12p�b�١�S�����d�jG�Ys��ϷG(��ڍL:�oo]��Y��c;�w�WP%�)�?K{�T}��������學0z=I�6��o�P��l+.��ɀdh�{���2�����=%A�"��%�
0������j&����r�ҩ�(���?�����n�J0�q��V-���-6Nӆ��^9��`�o���m�ZKM����I�a߭4�ϲ�+�f0d$�	W��SP�c�5:�c�0f$���,�k��Z�V\�y��읆p����W�����z��0cSB�k����xBB �����'����(�GMA~b ��g_�&[��8�������H���^TD��y�tS�Q�s,\�1�6�nQ�kg?f�qOѱ���-��F��
iR�Yg�"��%d��m��@t\�v�lnh {�y)+���E,���Z��;�~�w��M(գ�i��鲚��E�*鍂$�Π6��9����s����v屷r��1x�R�(�R���nZH
�^Z!x� �Z����W�('�/��r)[��n�ۄ,)����^y�j76��x�^}}_�_B�E��>}@�ب�f|,�	���_�ϰ�ۅG�#�6$�(�Ev�������Y�E�~�j�s�l��][Nv�n��G�/߫E\]�)y��~Q��d^智m�S[�U�o���������pW�WȺv��-v3� �XW��rzKdE�'��c-�HtH5�Hw.�/r� ���T�!n@7��ް�hs2)@��K��(��Pf����O��+4�;Qo
�(�G-�������nӚ��m�U~�>0*-¿������D�ym��ph[����M��󦹵 ��Lv�;8��p���۽������!o���f���ҫ���c\Z�A����h��
��_R*\;w�����;�/N�B�x��ri�4(O��^�W�g�-z�3�fH�X$�Eٌ��yg79s��ӱm�UM�Oc�6�Ɨw�,�]1bh`WR+�Ƙ��c�]��ο������d9��Qh�34��Ȟ�>���bC�=B�+�-�f(n�D��V���+m(3>� s�:��=�������:x }Ñ�I�}�W��/�/���_�����6V�ur�twJl��+�!bN`��M�c9m�dI[���}��_mQ���%Lǋ���~�_�4�:=�������Oo��p��V�+T`��S4��n4Þ��x��^9>Ǽ|4�*(�#\Gw���q^�"��9���M�8��6�����؉Ij !��ʌ���D�a]���!	�ر�J`0�ʖ�fˮn~C�P�j����Z���y��qA[��1}s�C�/?ǁ@��Ĩ|I�y҅_\7?a�CX��#S��m(��'
��y��~�?��8�h׋��0=H�f��@����1����Ex�J�>p��'v�n6���T�+��)wA톗�����������h��99�B�ԬW~/�:�e�G��i6Ue�<��U�6���'ڂ�j!��! "�W�D.�� b<��RY ���Elŗϛ�֟�T7,��LB��eN���r(��x_���Z�~-��%��Zw#�K�,�Zl$�i@ip|�e2��_��	��+���J뫉�*��K�Z���}:�E%Ǡ���=�9o��A���zۼ8F��o��%���N2�)�7˒�F��*�����|KAj�uV��`��n��!�O'|ٿ�^��V�n��+]f�n�n�~X����N^]� �}i$Pԫ
����B�6��PŴBzd���`�:�[H�/?� �poLP��B���E�m��|�ϼRT9E~�_�	��o<a�B��D�ԛ3��v)����ڵ��9nN�&�4�o�:��s���.�
H'KQ�-�y�?CNX�n�=Q�c.ȚK�8˴�y���*8b������j�ҷou3p���vN��
��6߾h�:�5��h�D�1�d6�C���$l׺)1ŸF��%�h0.>�
{��L6	���\��hr��B����13�ߢ�AI<�ұ����ϰ��2K������&��y��g|����ǥ�`�BFP?�C�u��AL"S7lp��B��m���mcJa{��ry?�)>��A�7Bf�M�����ODӮ��w�ڨ���B���7`ݘ4:I�l8#̐���5k���y�샅������"��$�PO�$� ����~Y��f!���cp�4ԋ{�*�������F�J�0dp#�pF�1/:�:�J-�z��%n�|�ի�-HXTa�K��g�_�]�x��e4�S0���5�����ˠW��:�����)1���_�]O��2	0Z�c!�;�Qq��)���9�l8Rk��|�-��>{�9깎4�^T�v֙�\�	����wmu>�y��c"��m������t�/h�{}]�Qx���)��G����H�@zU�n�u^����u(���[]Z����ɎǙ$d�Т��k�<��W)�����ܹ٣&2J���j������>�����7�:T�Js�C��C���5S�7��x@�U���R���7���^A�N��|������+'H[��S>$�'����s֋�d���-�1+�_P��~vk��&���soz���2Ρ����!sm�A���[�����w�����w��A���t�af-�E�O�l�}��Z�F�����M[��8m��J�"�܁��:�r؉j�'^��t-��R���`��'L�lk�:]��:�����4 ɩ$E�/��dZa�3/����'>�$��C�d_D�I���)>j���d�A���X�)rV�J�a�6���:I�����8��+�-X�r�9�I�qz�������a6�tDh�J#ab*2���2/�ٺ��5�nH��)%0��d�ĩ#�7`��AsT�q�b�G��u��3�3��ĤΔ��)aG$;9�5)����_�/�V�d�K�;����u�؏yPh*�:��:xl��ok�y�l^`UT-�Hԫ$��Sy}�n�)����I�K�Rn��+G8'�Z锆�	�	���[fS�墾c$XBz�l�,�`���O)�Kd8u.G� �0I��U���@�Xx����01�b=�̆��2E�ѳ�{?}��΁�7ϧ��;Շr �WԡU8Iyo�5�

��(&�ș�U��Z�:=����2�u��O�;�v�&�.';I�6��]m�]�M��]!X�ؕ�"G�]̳ߤe�w-m"�蓗�c��ؿ�Jvo�[ﱏ�Ǩ�mB�F���!
������}o��J�,*�*g)�ʹ�_�f>�B���N����(����ؾ��_2����V��ha���i[��$��or{�x� �Ⱡ���a��hA-��m����R-
�����<N�˘�\�`K����Q<��Y�H2 �9�0OL�gPxh����K��KO��J�9��7���[��9�SP*��=#��Q>�������Iy��wo�,pw��aܼ��=��a`*zZ;�����N\��9GN�>��8f��;�^C2ߞ��_L'��G]7w�{��r/M�[���R�$�.i� UP�lX������7t�1�Ѭ�v�u�]#aRl�]1��:L0�ա��V7���#(wp6�bH�J���][!kI ���%�ED�H��݈�y��f֥칆V���w��ľe�r�Y#wa'	d��en-�s���)oq��K�J�Xa�#��L�����81���+�Yʣ�k�$���N1�� XS�s\�~�a���YfkKPa/��.���1�����H�[���م�����x��;��P�hpg��#'(�5���?ڽLp���X�_"�&����0s�D�������H�k�"U��`���΢ѩ��c�8��_�a��x�Ҏ�8��¾��������.5��(�eac�q"��X�`猿O���*o(�#��i&���Z�܉��/������ \�:��<7Ԕ��.Tz[�0�R� �YG�b�G�V�DT��'��Z2�(̕� ���{���5�`<��͑�H�A�7t�n���D�I������
��s'{���H�S$�?w�X+g+1�	�,����V�b�x�@�vg���ˊtC�W��������?	L��8��4_7��8��)M���AS���M@���<.�e-��^3�V�����;���#�}�X^�Y�����Rb�{w�6O����g�{ޮsb8Z	�xg�/(�)Y��!9Gk�����#~��`yj{�?�bg�)ha!WR��e��2��9��H�Y�.B�h�!�����͔(������`�����6�> _�%��v�k���&�����DP��߬�q�w����";�����)	�����~])����u�↿a���j���AO��Mڿ�H|=�5zoUe���oD��q� if��k,�*�3�H�N�������LJX&�������-0�^M�l����JK�^]�x����2�C��H(�]����ᵛ΢N!6�?0�u�;@o����O�XBo=�e�K����[C`�,���N ��z����da�>��QP�>���J��A����HBk����?�03/ЏD����8�W��ED�#���ĤK{��-�|,���?������J�-��%���?�o��uGӧ��Ȩ�ǯ��1�����ˆ}8B�,���ӕм�c�it�J{E����7Y/��nր\�?�SlHf�H��q��LOdy0����'�mP�a1~	&J�y�?����̜�}��be,��j=-ݼ��"��I�#�����0�. ��Uʐ�K��Mz��:9Zb�N��8'Y�܁/R��G��+?a�D�����K���{�*e�`�<!�&M����iL=U=�*��ՂGr�q[�]�G(D��f;���4t����*e�*��;q揁D%	��C��uYv���V�l���Kd�����z6��k�h<�α���qE)�Z_��q徙h+$ڊ�u��
��]<�� ;!��"1� �����6��P��ɞ�/H}8�w�2��F�y���fvܧ[�9f.��(NT�|�j��~F!�B;�s���r�'�g�O(�֓��jz�����k�to5�=9t��i��vN\6I{{��6��i+���Oe�����9�ӽ�h��J�#�n��U=���&��:ty��n��.�<�{�}�b�r �MC��&�����6ZCa��{����:b�����0�T/��1�l�¦����)g�]Xē_"�J~!)��v�I���No��˯n���ΰ'������OEM�� j�ї�s(��v�����j��J��*�u|R��1ڟB']����}:���%�}���3J�u:y^�0�J}��$I�����`�!U�P�d�"�t�*�h�A�2X
	��C�\��ڡ�\�=�����Z�ҡ�q�mn9�����urňr&Yp��H�wGO���&6{�k�˔����.���5�L	��Ij�6���Gm��c�*J�o;���֛?:��}��c��ݞgs㶷�݇}!����N���3����#����������X$ϣ�����K��]�湺�ߞLѿ����|ƹ���%�b�������%I;(��
��\�u����X-��e]��%Ǹ��F�⛉o6�|�}l c^m���h�rT9�V�K���a�m���4Ց�,�oeEW�3o�gc���J27߹PW|ډ��ߣ]�;lNp�v��Hie�Fy?l-�Q��� ����	����mvչr3>�a�����2��`5�3�,U��1w}W�]+�RT�_5W'��W�����$�� ��Zh��l�v����S�|me�D:|S�)�kX܀l�h���VKƦ\�7���w�l�:6�X��Ab?�ʤ8����-��^BD�.Dv���O��J9v�"�"!4�#�jU�Dtv�V[������l
܎�J�u��|q���HW�ƅר�y��֜���q��t�9k�`�F�o�5 �$n��ر:SA�m|����\����A��ݙ�i��]$�8��(��27�R�2Zz_f���Q��f#���?T�J�,�m�f�~�f���#���%�e��J���������ČzmVxe�o�"{�R�K�^�p��fg���KGo5�33Kj֩��T'Q=�һ4Xj6Z�X�a���]�;���m�T��SD4���������o�3t���|��gQ-�`ib��Oɓ��i�w�!�=tT��ފ�K	 a�ۘ	\��Y&���SL��k�b��h��J5Th�7[�a>9H��*�t#��|�_4d_g5���%QM������φ�!UI
2W���D�(���Ю�{�3�t������3�%%^T����������t���'�jܪ^�y�W%h��>s@}[@"�{8h�'���V]d�S��mͥ����Z�#H��^��nG(u�� �}�9�`d��#ܾZ|7����\�!CG!����}��>F[
�Z�T�$�M�`�3����Coo�i������ѤT�~��y���P�k[�#/��� �Uz��]ҧ6��&j=�ߚ���Z��_7�B�Lc���U�7xo���ۨ�k��ӎ]V�i��w�n`�h
�kE��O�澬�k|+�I��YG"�|"'�F��,$��3Gh�:��-��Nr��cZv��q����M��C�Ʃ�˘�ʼ��=�]A�ǰ;�g��q�+RdF�sx�5�꒩��,+�eo�S�<O�+��<+����5�T�<z>�&Y��*q|Ғu���s��imq7��ZoQ0 h�GW@�JG� "r܏�V�è�ٵ#�\9�f
"j����s���a ��+�@�!K7Z�S8�����W2��yȄ�HP��-t����]��ܻxdgstnp�?w�u ��FM+2c���E2�]T�U�����wI/i��&L��yKip�!�&Q�{s,���9�'P�*�����������JaT��=t��?���0��}2r4��S7�}�T����k^�{\��Cry��堩l�H�З�F?��d���Ɩ� ��`Y�5��սgr>�1���^�����Zp�)�1�g��W��'����W���%��{�njl��-����0��v�Ê$�|m#U��UE�ػb継#��'��_Q0��4|eT\M�-� ��L���������w����0���ww�3��Z�יuz��K����9��8�y�O���v���כ��K�s��]����تh7$rP��N;�L�׃O��S���
��Ϫ\�96�}2�\v��MR��P\���ݷ�=�=�]���Jz��(
>y���.Q���.�'c�Wg�i�h�S�� �t=����-^�P:+{}����HYB�.�6�������DT-��o�|M<��`��o��̷VԻ�������OO'V��6��HU���&h��>׽'b��)AJ��938nY�<�b<��N���8�[+������Gx��놮��FWL���<�)&V>k(���mh��_/ f�����;����}2�C/;���au(5BAVs��m���ꍈ��~�I󞰹lb�5۳���'<w�g����m�If̉����3,������'�<k
h�uZ���0�����V��������]o债�;mC�-�`��� ���&PY�J���,�Ͻ8@��'����4�7����w�sl� ���g��:`�-����:�]i����7k�k. ^���G`�W��y]@`%���uLX� P ��	�4Ce��û�!类�H�f7Av� v1z*��WN���v�`+��y�* ��6�^f�,"�#h.��ǰ?WP����&�v�^����2�����͓c<���d�_I��������Q��bEKkv�*�/�<n�(s�l�e����wT�h�^T��������$�}���I2����zf�ksg:6dL�-X��;<ld�{��s����e���j��	��q���n��O�%����8��ܡ�䝈� S9z�8���ô��2� }���
*V˵"o�ыr�2��_º**�]2k���8�D�v]<�����F����+���{�U�V(�	�6����8A�A�r�]��n37�PG"�h�!�8��ݸ��y��� ["�?w��@Zթ�ʟ*�5���� ^z����g���C�t������)��G�$�e����Y�ev-]yK��H�͉�����&XkW��WՎ��`Dg$��^OW�H)3տq��=�.�K�qO��09	M��c\N��`0��TL$�K�T���\������&��r?���x9YM���44�biG�:ۦz���x�D��!~0�Q��Vo�7����`��l�+oӭ�R;���AH̳2=F��ШD;�hx���#��ۼnlM(r��ނ�
3���a�����Zn�����^���O��|��}L�h�Z5:�JJ? �-��d� �B�����ê���N���}���n��m{j(�8)}cGYP-�J:e2H?6v�T�W�G�&n�m��ya�V�@��Ǆ�$�S\0�ܹ
��<X�8?|�"�
n����NOZ�<��u��F�9�?#E�����O���"�K��`�)�%��e���@�#��~��I2eԤ:1�T����к��j��c5��֧�x��N�8)g�(^0 @�I.o��jғѴR�fx���u��QSu�~�5e�n�������e�*C������k+��P)/�9��K0�����P

�e�&x<q�7���a���O����G��Җ��#._ٿ�07v����� �ώ���gA����YU�ߧZ�K.��D�Xg6S�L��k��s8��|�N�D��C�~Q<o��9��^|C�G-��UʆW��m��J�Qsɱ�¥�~�m������+{8�����0s��[^g�I2W�e��<kFv�L�ڒ��5�n�^�*�.�P]���������/��<�_�{�C��;��U{n�h�?˒�dn��R	s< ����8:^�C��Y�h�7�=$���Ӂ���	�ڰ$���:�-}�jJ�c2��^Z��)�V�4�C�\g9��79�]�=��q�|��������։0��S��䩮	��J|,t����8�J:��A���aD+vvZӝ��kH���_;��ӟ%�M9
D5��嗑jQnk�퓄5�2��I�.	�Eok�,]�C�Z�v��l�����( ��<���kBA�/��91<]����[ѩʌ��+(C���N'�&��%�%x����Jxn����3jp8>�4Oے+L����ߏA6�:U�%�SKwT�ב�M�>w�,@����b[
�&<�s�!W�����Q���M����j��g�g'r�@Y$��ď���[@��8�<W��W��ȝ�1i>�V��>�Z��\{�98�,νƹ[n�yd��HS�����4����GK��R�mR���]�=�<9��a���.'|kD*�>��)D2��f=����B$#�х���Ӗؐ�L���ׯ�Pԙ/�ȩ10��6W��Z��vC�0<�UX��x6z�C��h�JYf�\��/O��z�F���F���yĈY��"��'H���H������N���C3}��@��ibn�.����*]�MX	P���~�ʉ�kj�R��z��E��A �Y:>>r�ɉh~���w�{�a����?*hO��/��8�w�`>�����z
#�ԝ�R]2je\/Si�KA0h[3��T�� �W��k�|���FG��a�����zS M�1���zJQ�+��̹"�z�%��M��0>3�\a�MY�����<���o^Ǒ^�gV/B�.h�s�=��<U��f|� y�0)�0�&��L���G32���RR«��Us������D�FL<���M�б�h�w0A-ҵ�[u�
gp�ļE��A�K�,dn2�C����Ne�j�5jG/H�T��Ԓ�r~��^� �|&�&���T��L����X-�\*��Z$q�iEMq�]q~R�N2�b���Fv$ _&�C�C�Tcy~�6�Ή�� T��� �X-�l��n�^��d��b������&�bg���GF��ݹ;t��	޾�xn��������`�_1���?"�\ؤv��dk��F��Ѧ�t���)�ł��yu�?�`̢����7k��Z�ň2"�~ʭ��j�h��z�_�]B,%�[���+6I��LK{��^vi�Z�)cvX�FP3��ֱ�=ଜ(k�l�g�:�L�h�i�ވ�	ʯ1���e�����]��4v����ᩩ%>.�!��܊
�z�����xL�o-C�.w�����~�����yR�T�݈ݏ����j�2[y��"��XU�Iܰh���ǰ��3͎�E���	��nL�g�4�+���y�6f����;���"好��)�|�~٩]0�ϸ��d�F�)6;�Y��*v�ഹ檧�c�y����}�cj{�}���(�g3�O�������+(+._�&��kfzگ��(��f�)�@-R���KLc�8��ߓ�w�6�}�LaR� �-+CEi���D���ͺj����W�Ga�5A�n`'g����"Ŋ�����V�W�Jr.R�B`H�|`*����涔ک�) �$g2��c*�?�H�kYY3��h,$�FP'N^K+2��4����z�Z�� ���Mo���f-�6\W� ��"��َ�X�Q�s]
p�3�� ۸ ���os;�np����Z��4��Y��'M��9�&Jjmz{�ʺ"R��>�'Y߬^*�����pK_.��+�fk�#S+�tlZ�̧SsվSb�2�{�ea������^��\���c}�c�@���Ӽ0,�S|, Oy~~��f��ֶ��}{{��w2薻�nNJqt�.�B�q����X+�E��%���9��y�6^)���y�D�6����Ԏ?^���k��	pƩ�s�����?��[��Nb�wRk�1��)��4ݻ;������M+�x
����_�UOu��@Ax�4߿M)M	%v�ޫ�qo%~�ݐ��s5�}�1���T�%���f�< pG�[P�ioo/���ܻ[�Ɔ����I�g����f-�t�9k�7	�n�k�^)5��F�fc;��!��u��1�Ic�//=��Sl���>Z�u�
�O�Y0-�p�=��Ɇ�#KZ� I�$m_��{��Q�cK(�m�!jwk-8���0�C��K�М�#����_5��7�a�7z��7>���8�l
،Z�Ch��M]&o�Уʶ�0��e:=rI���@mgp�i!�pE ����~��]`e�.Ƒ�EEM��r�D���*-mj6ȃ��o����,�ʡ������e>�j�e���jl������ԝ��*U6��&�)��Ө�d'���kb��Y�"p� �N���/,=)TXn����h��
ܼ*�ɝ���_i�Ͼ�f_vs ^�B1oL�C#����������4sED�<�m��N;
�p�l��ʳ%D�s/]���L�DJrIccrK����nIj���)&	^�E<$k�&a��J2,���p��]w�G�����	�D?N��m<��'cͷJ޲�<5�c�^�
a=��W��S�2/�oT�<|n	��x"J�i�n���Т�&fXG��P�}��5J=�2����h�vZ�0`"�gf�.-�a��	���}wW�~��������Q͊�+)�8����՞v7n��np�^|ķ#q����M ��%H���W� h� �9��ED�����R���W=)��>v�of �Q�w��s�umN�t��
S�r4�*#H3���Ԕ6.���J	���z�
sx���^�b��ܞ�d�Ew���]�����]]|+�$ҙP�p�NB�,��&ˣX��Ʋ���x�� c����肬��M/[����bfn.���S�<X�/�H��΃�T'�v�y���2�ۅ��c����t��#���7��w4���lx����T�ũ�28��;~��Z�E*IXU��Xy?�`��yP�����S`#�%��FK�hy��Z("ӽ�kvv��
�v�������
iX%="�|����5����z��g��/�M�K �e�#�"��Kc �B�x��S�e�gl���o�@Al�L�6{DO��]CH~£[��@���oz)J���m-�a���xT���*����T$'��d�e��4<_�F�m\V�K� �`:_<�Y��8ܘT�� �����|�r�f���i��$d�$[N�O#��7n:
���Q#�`t�s�xJ�	|��&�eX)�T�?3�dS�pk��8T�?�i�7����#�L>� 
�'�M�����Tr㲭�#�T�i�,l��Cȥ����-��]��:J�zU5��=q��/Z8�'].���ץRE�~������aꗙ!Pkrr3h�G�뿎�Lɖ(T���#�{Dj�w9����I�`�e+?x�u2s>;��F-Z�{�:��AʆStn���UUM�5N��%ieԹ�T�.�(��mGس�t?��>a2��t�1��������ɧ���	�ث0*�-�O�E��Hb���Ɖ$��eC`�]�H0w�$�Fܹ�1���ʼt��sФ������@����̜�=إ���57wn�>4rc�����o��}����w�J�1�Y���Pm���mZ�U��y�QW�ԃ���TN0�������N�� X�a�� �䪤x�q���⫹�~��1�ېu�7n�I�^�%���jW�d����dG2���M��W��zx�9�~�ajJ���B12�n)l#���dË�N(
��_�'b�T+	� s�:C�ҁ9�{�`��J��TN�Q��m�jc��Ρ2�NWε���h�����(�f�}N����Wp��⦷�"�m�km
|XÆq�M�,{.
�ɉ����`u�-��Tn���N1,%%�˚߲��H�]Ȗ��n W���v�*���K|�RӪ�y���ü`&?��-�2����䜁��i� I����'ѶKq�p�1��7a�j����I]ɪ��{����������o�ԞW��������챊��e ���=��V�{Gg�r�\t���a)/c3��_Z��4ҩ	]�|QL�v�T#�:*��W�kL��D� ���v�C`��c��ܧZQ����C(�r[������Zn�:I�+�t3�"Fׇ��a����B�L��6�F�5j�1�ŝ��@�d���ؔ�c�Mg	���s�ϑ�v_��H˒�ڌ~�
�Yq$$ڿ��^XXȶ~,�&��j98�d�m��&�hqh7Y��􍊑Og�B�1�E��5��f[􎢼!�u|:m��Un3��h�B���E���\�}�@��AѾײ��訠/p�5ŧ]۫'0@	����$��@
D���<�nfs~>�D��\���N�3��<��"	rXd��2��_a*�ws3��Ύ��ŀF,���͆&��s§I� q�OP��7 F��ݘ�;����7(�]+Jc�_Ó��u{�$���j�b�x�s�[:_��?m�UV�T�I��v�*��Q��2���<��ԇ����J
�4(�~R!�<Q�{�T�O�����b>�����;(u�v�O��f<������Z+b�3-\�:N�O"BD�c:D�ْ�;���:�G����{�=�j����=�7)7���::D���v�������Z(��:�xo 茏iY�՗T��9ǉ���T��ja�����l�TLM��V�sN(��장�������G��Ѓ�J8��l�NC�#$�V�&�N�_��Bͩ��>�ñ'�c� 9`x+M�pH3��)�m���a>��ѩV��#��c��d�}M����&��D�N��N��[���)?S�~�%��N%���i('/f�X9��3�H�\I�݄��K�\��{�[w�Ȁ�LY~gZ��o�
����!P��H�`��[���^��{\�iA���V�IM�n���Wv{H䓷��3��`��3$���i�υQ/uZ�X"'�S�(}�@��F/�L��Q��՛���8? -E�ZDx�^��>nԄ���>I�o�~�t���4�u{®x�΀9m M��5���܈̓�[�J���nnk�>{!�Õ���M��'7����ux�NW�7UF�绐���{��**�����k�b�B���jV>~�;����A*��T[���3>��#�G�B,�v����l�+",�p������x�PiGA��8l��N�߰�jW-�՞2�V�r�mz���RQ~"�AR�<�^i؏��\�Q"�,O0���%at�)�hY�9��y��p����.9�D�Zh�ځ�0��g+����Ř�u,e�<�!b﫥m�2�7�o���q]��#���1��i��b�mu�w���3�m��Ә���?��1�� )t�D�g-O<�|��2��B�'�	m��k�O���@H*�#�mW{�NB��0����Tڻ��ר=�$�}|����r����Y� ��\�������΁�\��l��5�ȼp_�2(t�J;xK\��a���#}7`��Q�%S�X��.���.i�w�H*�\����A{�zaF��d���-��T������5-��~� T�s�n�]v����%�V|���,_7+����ݣ�g�����$V�%���J4B �"v	�᝺�i���� ��ĵ�j3���^KIh���߁�|���W�S�&h#nkL�:��[����,�`��>w�>�R<�5jx)J!b`a��v�PiR�2]��r����)c^}��SE(C���_/4׉�w��M���#��[_�������¼�1�랟j��f��)
���y��T�8��e�T>�]��4O�r)��Т_Q<���"��4L�����)^b�L{-I)Chӯx2St��>EqC����	v-�g�+u����'���ot�������	r�s���+Z<i�iL|�PF�0ӵ.�i��P�y������C�B��B ��"/�Ы�3���Q���o��쩌"��Mf�?��2������I*��
�;�1�6D�[iسĪ/��J$��6\���&�ی�n��x<�R��ʭ��l��˳zװ��IY�`�5QE�kY*=<��.�V��$o0�1�x3'���g�.O'1WT��b�c�ZQZ]����|��'%4����� �jv�c�B�'�ُ*��� f]U�.|C���H�]�E5��@�[;u��Q�c4D�Â��qpTo���L�*̙���o�M�ۭ��aߟK��2���z�d�V�Q���$�9l��?���
0����,y>�G8��Ovs����e�Z��9������yv�X1���bQC� ]g����Y+V����ʃg��/s'�?w�)a[�VT�h��x�$,�t�t���?�Bf��6��l�jp�����F�k�:��M+��l��g�Y�?�Hq1�9x���6������&Ҿkh�����dP�������孍�W�,_�I��6�p�<��p�|aa��~���S�]���o��y��7��-q�(�rZ��-�>�M��!�\�� ��RJ��V�VZ�����d��?��:�$r!����T<,��5Ȭ����12�K-!HǭK��-��lݎ_}�׋8����0ִ��.�b��c��H=s�l�J��-|��<��t;�D��#_B�s�Ҥ��QrW�� �ɐ�K��ܮg�a�ىɯPת;Ͽ+����Az{Y��j�&���9K63��NC��jߌ���V�1��u
�Z<��F�rU��0�)��z�i�"O�>[�cǥ��g�C}׉�Xa�tvŅb��WF����o9��S����r`{�~�)#M'�-��8�"����^�i�YfI��7�9Kσ�AUΝ�&�ǋ`�z���(o7 R��<'�LQF�bb���+�ꋪ�����jG���)��[?p��֪�j	잴Tַ�9E[�kŇ�?����N|c/�����>���Ĕ��0���L9d�w���x]���D�գ��ȳ��WxT��n�a��}�y����M*,m�moT"t�����pu�u��u=��Ծ���-�e��oI"��o+.c{��d�|v�
�0c+�%�v�Y�jIZ��}�i�M\ߴEܱ�;r1��K�]'� ��q�c.�u����y�X�;6�f���yLR>��ഋEKo�(��G����UJ?�H�E�ſ_�q ^�f�]zŋL�)p=�C��嫻�=���!"!b����m�>��1Ҋ��]i
�X��r�c��˓�yA�jS��'�U�Z
��Y*!V��=���� ٨���.~/�k6�̰G�D�}�zR�� �:CU%�@n����&�C�f�K��HA�_��p�e.E	��6S��!���̸۝��O|w
�@��T�,ǡ}��r�&L$�<����؅g
��:�{ťsR�;�ܦ��o|�w��Ԕ����
&GS'H�-�Wڇ��&o~�8I۫��1�O
�*6�KG�,���m5�����K��as��Ջ�;J3��)�r;���Ʃ&�]R|���4J�TE ��i�'�i�M
�M��$�@�"����NO��(�m�����42	o�X�L]�i���v�{�\$�O6��lb�^��#"�y�e<�}Qx���+�Z��^|u�4|�$�{��S'�����@	��	yq�u��B�a=,�X1P�St�f�#����qy�%�_�w_�7 $x8X�x]���r$���X��j���S���UU�Hi�jA�RJ�X�U+�H��po�^L��^2=��<���WN�e�t�
κ�O�n�1V��6��G��T>(J�t���3ݰ_m��)��eΛ��8&5T��A{�ޢy�A���?�\���9�2�>�T�Y�v�0^������@���5��ܭS��ٗ�F��X�j������Ƴ����W�ݟ*�|:#���?������'�A,Q�uL�b�J<	�|zSRM#$���8�}a��qhޭER\:'�L��B���`6I���f ��I��zZ�9O�^�<���N)[���ק �C%���o�8B��$	�q���|����Y��b �f67�V�P��"��7�<�	X�@�Z(ڄ��)��#�^�W���`'��O.l���1��Q���� ��������t0�&�Zk��b s��"3����[�����̎�u'��$4�_�Qt��Ư���,u�M�9b�ؾb�DxH�t��6��1���{���2�-��DB1k)��H���r�`\��*�@�ꜫǝ�-"y����I5
d�I4X-F=Z,^��x���:�R���Ƀ��ޥg�0_Ec�;@�u2sn��Hb;z��Pʾ4_dښb7D��8	E��E&M_^��p�����-lu���Y�;��H"ؠQ1T�J3LQ6D� �Tzx�lu���U�Ev�����٣��\ӿ-�M��X�	�Z�]P��x���{�G$�y SL���w�[�_*|����~��Ao;cS�>�X��p߼�/�_���C�Zߎ��cV�Oze����n���X&`}?��ڻ''��k9�$�0W(���C�/K�h$2�t�b賃��imS�P�b�������$H9��#h�o&���)��^{��+��&����ߝ^@z��1-v�8�[U:��*Jz�Y�����ThL��Q��)��c����f��k@5�pZ� 2��T���{=䢯�s��?Ɏ���i_���HBB�`h��0E��R(>�-�phI�6�&W�siԶ|-�l:I#mfUȈ�:@�.�;�MH&���s@�x�����C�҆���Μ\��a�Y�U�Um]�I��<���X���W%�1�FC%zM�"H����s�p�Α�y�j�7�����W�ݗ�E�r�1��/l���*L�Vc����w��K���s�x鯗��L��]_�"{=������[����w��E�o[(eͅ��Ć��9�.Sq���ÜB$�:��J��p�v}�[JT�P8#�b8��M��p. �p�y��]�|�y�w����B�n҆yg�+ݓ��'�"�IGߏ��&V9H\M򹛻Mw>𫩁a����k��B�i��M'� Ҕ� f��ix������KjL;�nN�;��J~;�>����m�]�-�aX� t֏f�©�85�_���-V����������Y��bi�/�TC��Z���N)k~|�e����79A��n�]1�4���:j`�!Uw�����tv�}�b�{a�ngi+�c0����P���Z���1Ŋ�iS�7o���/�v��l����vS��*^V��ΦYv@���6�:�16!�I	���j��O_VȕWܞ�WԜ��3��I*�1� YG�%�@��蒘���N�qɞ�)s� }i\H��bF�x=�1�6"�H/*Ͳ�?����xP���p�SI=��HSo<�7�-�p!m�r1K�<n�v�$bEw<�Y�\��g	L�v^��YsfA�q�BZ�D>�:�CƩ2v25�%�^��LD=�h�g��O�c����u�m�k	�*�t�����)'O�Kmk�q�T)vQ�{FQ� ]�M��&!fI5��zS �WxxD�[����r0�ZlQ3q���j�B�w�o8$u�\�&6Z�b_�&�!I�������9S�큣Q��`>h/s�.�j���0����.���E2h_VfaH����f1m��'[�W���������,��P s�"B�_�1�J2F}���x9���M��1��9�)����@LL��m�n�H�.K�LAѣԖ�6����mC����2j��UE	�����a��!U���<1���er�������h�)euZ�=r�M3��|��N�m���E`آ�A�k�nL�Q3�_g��Q5���'��Q�2N��
Ҷ-�1�����v�����]5�P/�xq��@���:��79�"#銡"MrSզ\-ϳF>���__L��h	B�7ۃ�2ѓT3�*}��RG�%Y�4YU��C����t��~@&fUs�
D2�6�:f.;���G���=ݓ�2��`�Qo������D�������;��a�ZƁ��F�_#4_��!E������_o*q����zr6�}g����"5��"	\�|-�P`[z��ڲ	v>�%*�+�T��^STM�NF�#�K.�=mӲ�T{��3&ҳۨϗ�������f�z]n~]�j��pd\� i$��%{�!�C��%˨�Y��U�<z����Y�0d����ʒ&�z0�eq�ǿ2覨�vW� ��Ic��H|<��W.�|�%�b	��^I,0�D��d��&�{��k3#}(!�:Ց��:��A�Ƃ���ͤ�'AO�t���B�/�ұ%��+���uqjO�¢��Q7vф`�Y��"a]�RP�Gn^��"��l�+�WsY2�#M��m���``�J.Og��w_y�̷��q��i��[��M��!n�1�x]��L�����c�k?���M��A���p�#�Sd�H��Mڏ�C+�jV ��D��i�P�U��X����]u�G-����j1�r=Z_��R��}���$`3�B2��g��KjNנ/�0FKn��;�m۫�yGNfx�m �����}b��0�i��D(ڙ ��;"���ץ�=כyaG�',E�I�)�`K���z%�7I�]<���'K��/kg�?�TК��f�I�1�M$K��6�w�h7�&�.a�#�)�tX�e�쫽I!���ǜ����>�-0��Xb��J��Ч��ԉ:+?Uט����ge�C���N��g����:$7rS���e���ʹR����o�V[������ l�S�r�&��=��d�/�nu������/O;-C����S�D�˗\h��[�����QNT���Ά����$sC�DsQ4J��O���~>�[�_�S��r�rby��z|�免D~�Z+M֧�?�%��G��^1xv��A�z-�\A���2�?��{XA��lp4��2��/�#�r$⢺$|����M��N�D�������N �D�>g��� L|���������h�!LҸ��JFw3��/��(fVJ9[�����L�t4y��9և���k���G��}�iζbUg��T8%��e$.i���<�s��-�oLX6@0�,!� ׉���$�!�U�	�t�����Ӭc=Y��<n�w�D�̟��W
r�pQ���!��?1���ew̌�z��!g�j(&�m;�O��bF��scc�*�F��k����gM���9 a�B`����m�]��`$)~�A���P����-�b���l.��UF�i/IK�x�I�2I���r�[&�l%���(1��P,���4�# �h��~ޫY�Z������~B����RĹ���%X����y�R��Y�}��a�M�7cn&�gةP=ě'���_ %���8'����WO�����sk�W�M#��(K&�s���O�X��L$��0�#_D����5��A��:�����]��c�����8��& g����zAh���1��r:C6�L���F5�jx����\����̷S��	�J�	����5����r�7�~�K>j��|����$�A�W�w��[m��COT{�E��Bg�%�V�;͔�>�a-���X�1k1�K��S���d�)��]����<J��`�FV`f�pv��p���e���T�ePH�+�w��K'��l_�뉃�Z�� i�} ���I�����4I�$d��>e�ڂyi������&<`0|�H�l?�	ΏBYP�[�JЖ�o�V�Z�O�u����A��?+�i^���}���$JƱc4]�U�b����K����%�[��)W�x���l�zf.ۙ�x���X�\~PP&������AY�r~�d��	���E��v(��P�ߢ� S9!�T#�4�ЮC=��<��C�Cw����-��8ķ��JCF��ɸb��,��`ұm�ڥ���|*�����nT��_�uj0�$+���ޒէ������&����EV�-��*ڌ:tV��m �� �$�i�^̅?'�^�Ǡ��cHt�{5�S,>�9���.	S�߰��?���%�t�U:W�o]�F������Rt�� Ab���.�ԯG6�'Tn%���������D[���|�Gc�n�pvU�$��Ĳ���2��������������8��b�������^)Σ�u��.��S��	g=���U+T�(�l��=��>#��֭�%#&:�kwL����=ȳ<��M�[��:��|2�LM�h$]=M��e�2e���q���n�FCn��p�%x6+��%�?����������N��q����I
���:�qK���ɚC�u��u+f���eQ��ņ���� xz��q��|l�C4���hhU(������f�xM�k����3˲�~���VV&BRĻ����@������h��'ǕNN�n�.蠡J;v�/p�Զ�/U>۴�������n�s�j��m[�o���v�ma�7���t�t@�����	�-{�n�59��h�OC*�'���[��b5���p?^x5��Ҿ �� <D��f�7�}�!-F�AnS�^hnc�E7n�]'O�5:�a{��Ģ��C��B�yd�W)���*>�1{�֒�6"�Y5W2���7��.	v��ᬰ~��9tqr#3��o*��}�h��J����9wV�5QMŚ����r �<k9���lP�:�+㭣s(ʑ�jP��'��m�D#����n/e!\,�8on��Ӿ������vź(�BY�'��!�?nj�GI�Dُ�No.���0=m�$�����_C��)��9��ߢ�0:fX��ع�1���=|��B���0^=�9��ﺡ W\`]��d�R�_�׹��.2��vB���	�
v�8)��P�".l�rߪAH�v�M�a����~\LB�
f�!�le50����q�g�A�+�gv���<������ܽ^�tÁ&�}E/�f6��6�q���,D�l~��֫��j�K���~l��n������w�����wPON����7$��H�"�Q J�|��U��L\[o���1/�/%�Y���#%W�4E&��r� r�C,����wq�`�_-����{�HٻV��zI�K'��\�OO���ߎ�%|ܬ���y�;�64"����U�u���d��DJp��($i�Ϣ����6S窧P�;E=
����>��������O�"
���>AA��]��436����?��2V��G�+x��v�~��WV�d�oV�|�9李Rkӵb�p�Ϛ��6������ᄘ��8۸'q�=����p���Cx8(e9)�ѩ1s��~��v�U�I��7��1��m�.�����`�\?��-��y(�+�7��Ѷߌ���cˁv��!���Taˉv����y�s&��b�	���
ɛ���w�#������bA��ۭ)��r�٧��{g�i�eS��_����|���G~=�}��iv�v2�>��x�1��Uy��o� -��nP,����0��8��X�W��S���z��,'�MG��=�����߾:o�o��?'Z=�-��,�1��y���mn�\�-WK�����<�Ǌ?x��޿O�M�B�b-��L�X#ԏ�~��dB������'���V��j�r$

��e6`#��t�V���ԾlW�]��I%�d_N|&g�Z�=t����l��ԉ��hp {t,}���(3zXw9��Q�Ϋ���>L�r�F�ɵ
�ß�RB�hr��Uto����3j�����AI���xVXPa�Ngwe���?��~/}��Ұ���g�!~`7a�D�|ᰩ?Uހ�bȞ�?�:��G*Fj"Ӫ�bw���,^�P����j�u&�v�)�@���#���ٽ�eI$�	��/|�.�z�9�h-��5��3rL�֔���g#������\����8:'܅,ө
���~.A�
��h��b�k�9����U{�tvo,��j�ؚrq5ǩI��;v�aDؗ^��Qw���z�����|�O��y�:LS�"7�)'�ԵԨ^>���B��წ{�נA����kK+���ީl*�[�Z2Mҽ�=��ӭɫ��Rh�d\�S>z��S�ff|���1d���V	y��rJ�>�����x�s_�Ʃ�����qz�m+�l�O��¿.��ON���4�K��b�v�ˑ�n���K�R�B�?S���������PX7������n3��sW�`]�dX����ӱ`h�R<j�`�O�����L���à��c.��y�q�g���&���H`c�}?X��%�_8J�o�;�0�@!�!��Z:��������I� �3�a>��+�O��W���+4��89wG�I�)*5�N�$]���� ���?�|S8cރ����8d/��j��9c	�yV/x(������^�`)���d6�bz�E�o�r�j�2���_��Q:k%\�����)ե��3�	��lv�~�A5�%���nH��v�V�����"mǵ&�&7�޹}j���e=LO0��͜��a\���/�p�LI��f^i�!�ഝ�R�pJ��
A�#�ֳv�n^��o4������y���=��.��"LM�G��G���>������H�:���i;}y��q���v��;�g�4�f�)���r�T��,�^��6˫$|\נ��l�q�#��ئWcP9���O��V3��z���Ǟ
m��wJ�,#��^2dHR!���0Y���&\�p�F�l��VW1�X%���4��=}���������3�s�������6�L$��M�{	7��<g��Y��c}���Z*�*����N����#-e�����n�Ǖ���Q����Z.Ps�\l@����'Xs����Z℟l.��� Q<���L��64�8H�q�n��~6��rS����Q1(���P��I�鯌f9R���m�yU���'ʒ�^�:��<��}�p��*�@��UF���_ ��O����|�:$�`����Θ�� �(\�Uw�9���AeMv��j�g~��)�
#v�S`)&�x�-`^�j�՞�h�,�d��Ԥ#�U2��Z7v}Qǅ>E��̷؞�X�V���i���WrH
^�#]"��8x@��������}2"L'�+m�%͊*�^d�H���r5ù�6�骜��5H�¿..e��7���hq�c�\����.�w�t��(2�k^Ť�/d;���DN�֊��"�hn��v?��׶�|�:m��:�f��9t��M�~(ƃ#��'��1!�b��7�E�l]��x������^��	�/z�i��,t���!c��y
|�'9��!���z{" m[Kc�{47�ɸ�I��U��~�B^�Y����I�~�\�)v�@]e�J�ꮃT<9U��X7B���MQ�ڙ9�N21p���/��7@p���4�u��JN�h��1|�~�ԪX�DO��x�N�A�T���l�-s~-�5�sH��T��\TќY${q��9E���E����#4�b)�P��N]KnIٮ��X�^�&��@k����g��ly�q��KYaHN}�}*$�Q�n����G�n�\u�`f)�K?�\�?:7��w�=����G3��KH�~�O�*�S�;��r���c@x��)J�jl���Jߡ������Н.Д��X�:�~�r`Zp��f�/��$D+��������CZ\��w��9Fr���ԽKش�?���KA��jq�RuFn��
-��]yn����'-3 i$����X�-$����e,,�Td��^�Ὧ�բg�2�K��`;�Zb�9��S����������YB�������$Q79wi[�^$��5��4�\�1+*���?b?��)E,ߥ%�S(��_bV��|�B[6�h�\���;�@;�ތSk/(Z���� Pݳc	$�n�T��+��A���N�s�MmKk��j,���F���A3�V悂����y]�7����g늦��Lv�ߚ��	��̍ԩ�@��\C����6x^.�m���b]:b-;|��Wb֪#Az��0P4����֫�vUp%6�y��Ҫo�d��Z����Ό񠳕A{���{ğmMֲًp�> *fs���]�?��ȓXC{=ҍO���ډ5�W/�\�-.���B�wڻt�����K-l���A|]]�1�R�4�Qf�`�����^�k�R;'�b�/Qg��B��P�y9}Ռ�U�8|��ƒ��!O���XN�mo:Z }ܶ�'��Xùhe=�]9���v��!��G�*Q~�/?1{��d5��^ߊ~-q.T��� ��v��^I%By�؉h��Ew���C���^��`�[��.;��
���Η"��2G�#�3w�����uK�� s6۱w�u��t{v߽�_Xɜw�����۫2�����tP"<]��/V7�� �����n`n)>�0Ƨ\�Zoq���G6{6P�Uc��0�H\u٩�+���6�p4BḠ���q����PG�����o}3���*#Hsߣ��ӖG�s~�E3^=q~�k�Kz�����0�ҘC[��ra��� rs^��-�H�o,c]�U�����Ƙn`�| Q 51�[��{H����Ko����
w���Z�+#[RX�C����1��uJ�;���Su����c;�^ 3�������8;�?\�{��\���δ�����Jf���eu���n�.QuG��D޶��˖��3®���a�{��ԾtL��J����
���z�_¯R���ӽqb����m��@�'�[��� j�_uE����-��B���l��;�5a1�$p���`ݻ��ȧ�dX
�4&g���_k������ظ3�z�d��w���j'd�"S8��a�f����Va��c֍R��������L�&��?�^�A��Q����u�}�p��-|�8fJ��?�<�̛�))"� ���P����v(í�zF1��v����h�w��j�{F�>�H<{odX0�*�����L�~zb�04�R��B�xs���2+~�C��ٸ�ٸڇF��\��'8�E�o���Gw���ץ#�L�bv���<���/�u&�\���B//��{#��Wk��N��U�H��Mb��ɨA����G~�/�4�!�U�W��3��Rz��̺訩3\;�t.����r�ry�t�N��!2WC��]�l�Z��a�n�jј�S n��Q��ݺ��~V�Uhs�Ĕ��F�I3v��X�~�nVu�(�_ F셄�I�������B�j�k��wgM�����:>o��W����'DdU��M�����S1jw�3�9-1;-�Mf{��8�v�cԪ�M�^�_��\Dg��D�a�!��+Dz! �c�L�Ѧ��Gmv�ᇠ�|��>+x�U	�?z���S�//ص\�׫��FIfS{=E�_�n���Xb�GG�N4�rka��uU>iE/[���A��9�z=!|d�8F�xd�n��9�9l���ۧ��]b/VPs�iӈ-!�ᱵ��kH���a�Β��.x�����
�N�x28j�VF�ב.ro�@7��������S�ը9�4F�?I<�zm�=�"ボ�g�H�5hN�d���m%�ݫ�p�	o<��sn���D1|O)�<��e.�K�$��o��/��C%��!M�	,��1����-��Y˹>�V����Ok�NO�E�4�䲂���(>�I,��ʧ$����E�_o~}��d_HT-��l$y�,:�;C#s��ҳM="�-1Fι'�ᷬ7�LW�!O����~���gƩ���l<39!��	�ڗ�Z�)�j_X���0&��z�,7��-i|>�ܓ`�ZL�ո�!�����5j��:+ZΘJYp]V��o�Jyx��1'�.f/�]�?|��Sy=r�K��-l����xZ䖭�v�^d�+(]]/m��tQW?P��;
��K�|��r��"=��GIp����q�W�'O]8.kX�.&���ewt�6�*$0Ю�w# � -���̾�� �k������<�� )�W�a��3�~:�3����-*ymo��:g0jz��k�4Z�g-�.Gzn[mU-i.k��Y�]n���W6Y����
	���O4~'RN�LW�� ���\�ǧ��"j��d(c��9*���PM:e��瀎y�߂C�U?�OSݳ9hA.�4��!_�1p��g�-"�܄baw���}-:s��i�Ml��E���Pʰ���~���qn�	�)���&����+y%F��ᄸW�'5bP�M�T��uyB\�����]����V��#4��9�YM�uhq�9�#8.��cȂ���&�g0?�_�*(�+[{{D�o�>�4I�\u#ĭ���SY��Gۙ��k�g�`���{P{?4�_�kq�bg~㋱���g�6���%��~ւtE���Ok��q/��9Tf�JBq�t�����τ�ѳ�,6����WjQ��.Z~�0R��r=��(F	����H�(c
��k4�幨K֣F��i��Tz S�4�__'��̂�������r�΂���(P\)��7�I23WpZ̾�_̤\�Yy�3�Δ�t���ف�+�.��w�b�H���t�q��7f�
�|��:5Q�%�y�z^<��`vd�%��� ���Jf��h�w��H_���>͓i�� ��e���8$�J?�f���H����R]ge�J�v�D��r�ύ`2��=Y���'\1���1 ,J��d�e�(VDTK���7�#��N�������)�[R/�nNh�sz�&k���w��j������A����>7<������a����*���\ˍ��o00&�)���_<u`��	�B��GO�pvOP/���JLgA!�p65����q��������%o+�>�{j�������PK   {c�X�l��A Ԥ /   images/670050b8-4f2c-4603-900e-28b8075f4ca8.png�y8�k�7~��]	��%KE�N������C�Ⱦ�R�ꤐ=YZ���Rq�P��/��/�ݘ�����8�������/�u�j���z��g��Z��2�1 Xگ�� X���+�=j���U���� ��G��ϓ:��uW���cs��9�����I�OkK{�s��m��"��� � �W9�9�"ul�Y.�Ov�V�Z�d$�ί*H:�y���Ե;�_o�њ���>ض���)s{��c?�������?�#?^ia� ��Y[[��/ﮫ�ŵFFFÞD�L��gF�O�w���}I{�^�w��+���v�^3�Rj��o �зov{�������ϴG�&���*��z���E�]?N�z�Ff[2�3�͂\�$Y�\�p��v��NL�
�U�aT��?i0�&��}`���յ)��Dt�� GGG�Ș_�ҭ���y�8�X_U�hʫl?�7Bt�$�Mр�o���)+�2����G?4����%G�s�
'򟌌��?98Z�	zÆWt�	�����kk�s�r������J�ok����v�v�G6{9�ى�Ze�Vf�ޭ'��F�L�����hϴn�O����2S�'i&ȣG���"�(�i�4�"��9;�����R��Ӏ-��~�],BEF�̔�X�X��H`����Ư���{j�-ó��5
OW|]���YH����dm�j�~��uW�Y�Ke���x@�
.̒��Ʈ�����&f�&��Y����{��'F
�R����Gq�۷o�V����IƓ�Ñ��2~��b�y�D�F
�Z񚠃�UVK�&(v�_���~�M�7��~�M�7��~�M�7����0�y1��?�v�$�g�+��[�r�������D�=��DlM�ph֒H���\�����+xJ���?j���ܼὓ��?8�*D�I��x}�eT�ī�~y'Wk����H��}���G[Z�?1�7��o �fZ�/yQ��/�~���_����������T���0!ʩm�}�gf�a��R�k��ƍE���]R�)���Q �i�K� ��]o�+�+x
a&���Z��^�4X]���1d�*-Ԍ�ʳK�h7���Qu
�mKdLIG�("|�n�sj�����R��~�9[)ܞ辟��?_�-tx��e?�t?a�]�ȉD�a)� x�`�K��S��'�������1Kl�|�����aHnj� (�I����dN�g�}�R�U�e��{���?B>��м���zJ���2�g��Ϥ��!�B���sfU���Ś�c�x�����C��]kH��!���G;F\�@�Ȇa���\���{o��++{�,�C�R;I�[Ӊ��2�y��b�N��L�/�J���άV�^[Jzs����f�+y��>Ȓ�m������/m/��WFF����1��'pU)L��f�U�SJ�bH�e �NM�w��U<":��D����"!)K�.e��S0�d�-�EBD$!䋩�ܙ��H�1�e�3�� Ğ�����T-�݁��ޅ����֞�Jߎ �����!&Bk��R����qШ�9�*vU54���k�F�+!�4�A�Wv%*}N2$h�^WY ��E��e��Iņ��i����îb:]hNJ)�-��G�g[H��g @�'ݽ{�8裇&?S���V��̸1�@J�e�R�4v!XBt��1���4/ba�c��P�_q�8��J�ӡ֢t�M��`�����J{'�荘 ?�; &�OW[K /Q[	�pw��Z��Qi]���>k|�->��q��Er�| Џ�I@,��5Dn�IêI������"����e*򊮘(��>\�L+of$�M�2U�儐6g�@��t� �o{�*� ���X�W)�.�'l�GA鐪-��1bO;��`�I>��&?��,F�w������ߐȤ.�F��!*V��t0�L��|)�q�`� k>�'xM;�h�� F���q�Z�n_�����)H�+�v!ZOr8�7���	e^�4^��:k=]B�77�a2�j�_e ��/���+��[�x���51��-�.=�{6~I�(r)�,
�+vv��(E|�,�Ξo�^7;��QqQ�P���2?�]/9ޥ�[]ʗO�˼s:Eq�!�t3j����I���G�Κ�M�P ����O�cn~<65�*0R0e�?��6F�a'�[/�g؁���<�4��3��1
.S�N%�B^�*%"Ih�$��%ݶ;G��&��=��T��V��q�Kz߸Rav�٤���F3�%O�֒�/���K+��I�+���[s'T5��D�0s��QKc &�ۃoi�z4�Z�5���&�a��He���MQ�QF<a\{>��n��F�]���os�їbƿɗ'���?�e���t"�"�aAP$�H���6�ᢍ_�0#�2a�k�'��V0fm���	l���	�"c<��,�|���c�5%짞]	@���;�����k
��4,���1���z}���Lv6p����J��+M�5�C�E����NYJ���1et�r���7� Ds�خfO���Y��"���*hsq���/r��ɿ
&��b���o�H�W��5�����l��8 ��A2o�+��u�T���e�;p���b���|�zP͆h�Q1�d���w�y�I�?Vp_�i��^uV��EЁ&F[�A�fs���ҷՄ��oM����B7G� 4r��eZ�^%���?~��x���� Æ���a���φ��g�[C˜�5<�֭�F8�*w�/��nt����n��-n$�1�{Z{*�[�My��u|�K��*[��.��"�N�	�GBI��z�Ma0��t���).�u+�="���B1�d�ǬO��1��u����҉8P�(K���DV�Q����K�3�'vS,fpW`T��j�v���pފ�`CǙ��W�p�^���X�U_<��ƙZ�K4�*��l�CTe��\�
��WAJ�#�A������)-�6�"L{���}���F���M�0��`�d�j���pb	_�v�jI$�%�f��O�'��gmN��~鄦���~���fq�\�iħ�]؋.�o٠�aPT��\�� �d�������W���WV�X�mԽRz.S/'��m�(0~o��;ݟ1糖���9��SbdBH�iz��	��4�a���/q��5�c�@ ̾��CFkb��d�;��ix�aY�#�Y[�ji�ih�yC&���/���HH�q��'�a)�RV{��#�r�U�O����ceo��$�q딃$�6����l�8op��9�>�T�b�vI�������M�N���U�J:v-2�~%0����o�} P�Zt|��.�_:`���+��?����?�%� Vi���\�cz�k��\�K9=��9�a<�O���X�D�!3�ь����P6E��Z���xLo��&�a�C8ı�}{�J�@�`�4�)7��J��7k�e��%�ך	#-���`|0��6a7�׿F_�۪L���\�NN-\��#)��;6���H	���m����.�*��U�D�R�2��)�B$q%:�a��>�ХN������!�����d�{?R],���~1��	���Zv�k����Y1P�C�9�Ֆ2��^��`>��g1�<�Ki)�VC��c��px�p��5q�F��̽maJf�����x��\Z͖W#�����O�১;����A~�
��Q���l.�Z��̮���(�t��%�u�y%��2x���E��+My�'�����
����o�V`F4�ݹ�?� �(���XVd�]/rS�����ۧ�0x�#A�{2��J:r��~\y��_��.��X�ש/��I'�d��1��j�Hx�UVnZxV�?�Ue�b4�l@!O��z�?���C���3�B�g��p�'�T�Ӎ�y��o<�Ѹ�1��`9�q��|\��znQ�񯑦�Ƣ	v
��]��D=*�2a�C�x�[ͿGK��^qD����.�lױ�ֻ�����)J��|�QFy�_Qv��,��(��ϥ�H} �`H�(��th\���1B#�wV��0
<��:�nE�e��պE��0��ԭ[u����T⴬~�z;��9��c��K��$���u6#���?^��L��XO���O�JY39$z�r@�e��&�W7�+��]uV�UJ^���R����T¤�Wz�+����ldU����]�ݪtə�XѬT1���93G|�].0ʃ��jg���ү){K�=$�*��r?�G�k�ǒ����>�4��YÊ��4�JX� �$���rn�8��4K0���e'�͇d4�Ϡ��
b͐Y6����u�����/��0�i��?5�3� �oL��Z#�@~��q��l�T��Ɗ��Y��V�ϵ/��.�-ҿ���K2�Cɀ%����b�
�7���;���Dҁ^�P(��a�����sf�1��_M�,xH�
z��]�xl�� GJ)W�n���pkީ��EGC��?>>O��ű�J;�VW��w6u?��T�{��'��l9��_�{�Mn�6>�st!��,rȽ}��%����vb�G&��9���ʘ��7o`7�W�3[鰼QJ��Ӟ�!��q��GmLj�[r�]�8��H��H��� k&<��[)Ɛ^��M�?b�Co�;��e��=v�HWF��ŝ�V:Ac.z�x���J�]��|�1�;���K,%�,����6g�>$����x��y[{6�����t^D��ύ��6��
����A����U�'�6� ���.����n�wGb��ۉ5�xV:[�P�±�)u\�ݮ*�5{�[�%[	sdφ-여4D	r���g߅��*�OWKe�DCW�W5�`�)�ƴ��C��s�ó;�2�����Jp�㽻;���H���#N�t�: �����VZId�+�)U�H���k39�����"*##�X�Nh��`+6�i�/:��<8�y�-�$�CqyL��l�rl����o������X��^'����t7���e�����3��[	�F��r�p�U��3!�m�5���V ӱ��_�c�W쎬�*��7�c6��}yt2NHr�o܈�W 8��T�����N�\,��e�6��/�_����穥� ���E���6�| yY[�}��]%�y)�u�#/��`�)�r��U�W\�>lA��y}0���S���D�A�Lv �G�F	���u�J7�6�.�xm��l�\9��7D������O#�؍�����E�N#�i[i%��t��".Α��I�92	+�c=�!�C�0�Z��K�O���$m�����l|�r�G&#��ΣBt��	,Ƽ��1�./'f=g�^�i
�`�	@�a��hBQ��'����Ei�v��8fvM�<�"�s���3�Q̺�'~���O°Z�<��ԋS�
͙f�S[n]T]UTe���1SUU���h�W�3������o��gRpo�j�����<�{�[vb�9�%�^s�,����Lc'S�%�"cBA�v�%�49c�Cy�Μ�샏g�<45���1���
{�k��L淶G!Y)ݭ�8�m�3�nS�QS��3O+�m��*�0��9�{c�&��KJ��.2�H�܅�f�9-;sD���SB���tP�����{I���F3���t�P�),�����q��rT�Jw����~�$I���ْ8�?�b�d"��$)N<�3d�`��`�l�ia�w�ǅ��,�>K]�'�<
YX�0�;�j:4�A5���X���]�)�\�DeN��:���H�t�U��҂��<=���x�tz�}����hX G�ݠX�k���D�u�}o!w���Y�^����ʼ����d�+e:c�U蘣��F�2x�@f�(��m�^��EZ}ѥ�y�`atOX���Ң$����X8!�t�2�&l+D����28P|�f���s]ܹ�E�o[h�mY�@U*�߻�Zm.��5v���r�r`�	���9����9��2Zݷ_^ѣ{��lC��;c��c-��M��̗�.^4��e��ga�[��[��I9U<�eCd ȧ����G�;P3�?�f�}D��bb}'�h6���V�c��i�#�
e����3 6d�N���M?w��r����~����~�\���~��̒~��I����[����J�cѪ,�SѢN ��M��W'Y������"���@O�04^̼)#F|��	��\�'���*�d���f�p�b��da�bv��;j���-թV�� }X�N.P'�[?.�^'��#u*S�2���up�����q�Ξ'�����p���� BiT��R��"@*�����П����Ⱥ�YÓ|K��cA���,4 H�d���R���ێ�"��uq2C7>�����i�ԁ��p�)�t������+T�SKŗ���0�E���*?��,���[�z���_�m��!RB�,}�|Ϻ��<��F�}��l�2S2߬���GY��0��n�I��ʼ�>`d��g&_����n���g�brX������8t�`�p�R���V�o�L0Cë^�����-H�l�_�'�_ލ�,���xB;<r�\݂23�CW�~�z�s�K��潄�y�jŉd24&���Q�nȐJ�K���u{a�����g��xhc�����p�Ɔ��[<qn�C��T�����@M�r?n�:���&�{,�5oV1������[O�S2�	�E!�;fDX.�9���v�kh�ِ�ꛭ���g6t.үo5�U�ɻ���N�t��e�A
Y� ����:�*Է��qt�F`���{r0����HI����̄�V�/E�{;ȋBc"�I i�BԍrA}�[�������#����{[o�ԉMx�ÿ
��>�_V��E���V��}T���V
���eӰ�h�!�r8e�F�A+($m�� hN��B��U�W��(>B��x��E!�^��=��g��.-�F	h�r	���FY{A�.ǻp[���Ӽ�D�r}���������݃MM��ͷɛ��� -��'�,���z�u�Q�HMYZha�!kD>!�lI�#�U� H�5�i�8������	���o��Յ)�,hD6��Ɣ���q�� 7�K��k"w�����Nns�\U=��9�m�%�~Pn��7��[.���{#2���fr�G!��[��$ļ�v��1#i�{���/��< �Z 3y3epuj�uFn$W4��?�e֓8�:����&)�T�?uɗ*Ll*�����XG���?��T�ݼ;���b9?���塈���n/��)P�,���a��$��K`F�
�pJJ��)`w��PsL�,FQ�s��Q����#��co���J�o��px���vRe53�IԈ�W%T%����9��h@Gr��qDc��b-������aff� !����?$j8�%���xA����A�\�l���7V��ei�)͢��m�Π=��s��_�e�,�7��oQE��fV�q& al �"NND̦�=��6�<�3kzݓ�&dץ�|e�A���/��L}�t�
s��D��'�>��=1%��s���;��Y�J4�yD���6g�DF�}���J^<0��Y��t݈Ԉ��������O8p��CWi`�G©@y�v�%,���$�u�X�?cH����p
��� p��)�Y��\0�ߖ!�����3fo9fс�rH�}�" �>����Q�'�$�π	�5w�g[㰠x7���u��R"��%�/�m�q�gVK��[�B���(�)?/ ]��©�8�j/��$��2 �i�č�VF�����e����(�2�z���$���/���5�sٿ�ҥ� IC|(�^�?�l�������Ֆ �|#Z�����QGD�]Y�ls�Y�bp?NNY�?��� lފ���D!h��q#���^ |[�D"Dp�y��̼T�I=#l���M�X�6a�ƍ	��o�h��6CJw"��}�!���e��j���]��|�*�F�Kt{*tI�$O�oX}���3w��722��y�����o�{at���ϛ9Î�|�8�Cx��F�O�.l	�1�p��M�E��,��ӻJ�c�uu&���������fg�x��%� :��$o�x�����9Xa& ������;�yh��s��/:1��<�E�%{���_��eMn�w�'1 +-H�Y�KO�*c�xh�����M]��y�}N>V��8����\Hs� fq��>���>�,eee��[1�]�$��I3����pW���Sp^s��ٹ��s�Fj�,G�.h�L'T*L6UFi�r$�8�T�����<vB��bf*B۝�CKf�M�h��s��e'3e	(V�e&��J�|���2�/GI�/Gt!��Km��m�2��х8��z���sҊ$�n�0:\�zc�|���р+���g��*���:�f��43�\�Hܸ�`0�Scbη�|ĘE��0全�h����Ħ
g$Ұ#�R�[|F�9J�x��x��Gq�U���͆�YI�M�gj,]N������H�wT�?��P����Z�ј]�]1a|&>>�ݍ8�S���4z�۫���\(X��5Ki��z_�h��֋�s�����R����>�nz"�qFM�4����K���=�E=�J�o�@��?��{�Y�������l�t��fMnI�xû4�'!p^v�eϫX]�p��\��ff�h���w�oy����;ٔ�N?��y�k_񙹗�yH����q{�v�� �����\���B4�.so��|�#wދ�=�����˵��Zt�r S����3���uʥG\.м����p���hMr��I��ļ��αܻ���;\�A����.�$�q�z����b.�$��րd�*�Z�?i��$<���V1TWwv���M�m��/���O0���K੖�n2��|�U����_���k�XB�C���[���=tf3��C�l��t���:D� 8v@���z�SQ�3Y!�Px�ο
�w`�~`���N���J9�h���U��t��n]�p��m���sݞd�pd,�#���ݕ,U.�ߟ�>���$@sh<���T=3.{�o��@�I޴�g�h��SLc�ǣI�(z� ��VB��Á+���/k{.��І�j���.?uNa�=�3N�W��t���γţ�f]��f��hb5 W���ڜ�GH���xպ/��QM����)Tg���D!��&��\K*
�Qz���
m�yg��4�U��'�$\�6�iݓ����)wgC�K��;��{[�/�:m>Ro��GE�^����Ar�_�����Eu�V:����o؞ڸp 0K_�F��i��h���=(�S�,�[�u���E�W�X?��I�� T��ٔ��%���H�Z��,s>�����J��\�]��; �>�<
9f!;�8nv������N�Wu�!vr�}u�{�^��V���DC��^�ɯ?h*����B"��{Ty�h6[��^����Pa��1�<ym,?���ڌb���K���\JV8 OI�gVx�!v��b�H"����=�<u��j�"������]���5V�oh��My��ho%�B&H�~��:�$ʻ��`���q��~R���[C����n��ڂ�jP����	^��V�D�(b�M�}+�������2�F7������8Wfhr;�"'����۞�WR���Xh�QZ0A�r[{��t���1G?�!uv�}Y��: _i!��T�EB����t��ޘ�Eά��q��;�I(��[�t]��-T�L����S
^��[8�޼v�B/�,��7���?Y���B���	97�B8`��$A=�\)1��@�����+MJu[J]@�*��d}:P�P��^���V=���B&��54�n��M�[W�O[�'�V�g�Q�U���N��A�5^׷j���GԼ ��2�v�2�+��x��WvI�Z��2]�yJ-b��H��S���ș[�����ul���`^��е7����_��Ey�TC��&6���1s���EL�wo�D�tG�"�Y�r��k(�@�dd�p��1�o��=c<� D��]:E`f6J�k�)�QRqZ��Q)m��Ff�G\\rS���>G�!#��_�[�R�-��.m��/�:e�J�qs�`$QN4�_]�u����=ֺ>{UJg����bC���́��!�a^s߾�m��U��I��r+�E�s���O��ObHX�L��wr�H���!��R�^���`=0Ie˭{�KA���s��rb��W�)�6��<��`���8S�X�����ɔx�gY���"��a�')�X���J+F�V\B4�5�A�	Y��"Sχ��#豗`;�:QK
@��z_�kl0E`�MX����&?&��4r7qD�>�d�������> I9$�?�I�	����A��0+�K�����҃�qRL��`ՄoɆ)�� Ƀ�Nru��ky���8m��	��A)�ܑ��˥��!uR9�&  D��OM�q�tq��a:�8�a�B>�Tu�c,���`��ST:�T����ME%ϭ��銟!��ϋ�^�B��	/��y�ۮ&�-�a~ɷ4v�K}�Ur����:V��C�җ<�`� �I�j���P�;����Vw�߸�"+�����(�#�CH��	WV�}e����˭���X?���~��~��_`�P�3A�|���q�����r
P �����2�W�a�q�҅��en.�[wi����v�:Q�G�{�N��w:�H�%zF�T)�(9w����|dfff|Lt��T�T�n~v"#�`��"N_ܖj��M@4A�U�p�����d��Z�%��A<��)$($d\t��T�h��fG��s�����R��쀰��N L�<�>�J���w��X������C�}�3�9$�:��ۥL��:�-A��Q���!>�-Wi�j�e7�Ub��o��7�������}͢uan}*X�[R��{H�7ܥ�ԇ���\]gu�}��Vb��
6�����oz�'N�U������sH����7v���R	���8���͢	1.C�XO�'+�Vt�c�,{��q%~��{�.C}�j��*yB
E�
��0
��{�z��1qW�x�۷O;�{���-�d�.���Pe�����f�|nv�(�G�y��#� ��x�)� �k��	;� ���[SSS$3!¢!�8L	��� @��0�`LK�����yj�>'v`��9T��Ӻ�H�@���uv�܅��4>(�#��Vp��Z�*��\� 'K2��� ����W��I^�>�
4(���� �Ox���ЃD��>y�
���=��4�B^��C��(h-�Vv.�^������(wikd�2
����d�8Q�L����J��A��&<�������,~	?��Y����t؊&H�A�&r&o�v�4 ����H �?av囪�9��g4������H���H�.��a{Z�1Q��!4�ˏӴ���l��R���D���4��*a�+�>��]M3��6꤮��	s/c�lmR�m��n9��>�h^kck��l
L�/�@��́��f�$L8��.�r�~�X6��c,��:��<h'N�x��/0v��ܢ��L�<U��IU���#;h�M��ɉ98�͜�ҡ���U�QQ��I��ww�z=�SHq�">��}&pO��h��U����a̍�K�-/F����`B|G�QASk�� �*���s��A����Ș��M �bB!���h�����:�������\l��'��	���0ӑ��z1=�\|�x�4f?�6�	��HU�	5Cc6�5eZ��g�&f����Η��/dZ�[��t����"T3�t�'|���R�G��q=�{��ɼp�| 9j��(y']:��؉M��oC_�<,�D��.��<��*�K��6󫌳��:����p��1WC��k �ҭ�XPa�3�0�ј�'�C�F��A8ȚIx4�.4��5[���Bۿ3�r��qG��s�1{H�C4��?�L��oӷ�:�4h���z������������;w^Г{A�R��#�Z	��s��kj��+���l�q1��t 7q8vE,��V�(�Rl���b��Q2��K�ǿ�架]��0�4����l�r�:��j�^Pf��c�=Q ��ΜK�p�_�5���A�2�Rl������D"����GϮ�&u�&��Q]4�BB���Ք7��ڏs`��!V�a�&Ѝ��{��;~�=|5�|��d5��<�����L�x�W�5^���>�L�)e�;G�	�h//�wy�Ш�
��O쉾��ʙ���^���3�o�aT��z�rM�d��s�,��hdE�����?�է�Z�#�n"WJI_o�1*Z�3�f�q|m��-O���^z�G��oJ^��D��꼺�wT7Rt
3_[6�GC!�N��VuH's�׈Dq:2�u�H�}P�x��ڽ�g���1�A�4D���t�o��qΈ�p0��F�#������l*��3g8h�kC�2yK[X��Dm�T�{�x�V�O��{�Ֆ���GaM|$Q�M�A�rL:��
�%! ���{9ƪR�[���,�|ӟ��XN�&�><#%p�����,�	��5y�oW���nt�/Tێ���]1��z�Ldyv�1��lja�D��q�
��b��Z��|N�0��,�qe��BL�jЀs�ۺ�-�"��R��A�W![� �q�Ar}����x��:=ݱ�W��h���O�D/��ѡm�
��R6��vX��mˠ	�FB㞀�۲�dh^L�����-�����j�t$"f,�%��.Zr��ZH��ֿ�U�+���,@��^��4�H>�˭G����"=pY�m��b�,�(\��,2��f�u��)�S����ƺMٻp�a\-�*ք�<�ů�����I%{����b�-4�n��2�{ ����P9��y�������M\^*d����ɉ��!$�������p�����rك�R��Ә܅V|M5̎�#Ǳi�R��!�����g��~8�W<~.�x<	�>�;�/��k=h��ভ��!1o���=G�C�	���2��ˍ��/���c+���9j#�����:N�i%�+d{O��r��Vy
�=�VGV*ɣ�Q��SZIFD�1�2y��M���:�� �ᾦG>�|� �'�M�']���U
������K�:1�FY&'z-��*3������0�9���-��� J�;ixQ���oM%%nF�� �}E�/�L?
�,Mo"q�u�r�u�X�(��qS	�dH�"��n���q�������ST;���AU�0q���:V��P�"кb�C�}p5���h���X]D"�!T��7��5�i����{C!T�zQ�*��<B�|�$\ѝԞe]�MY�ӘG P/_�:
�#Z�Z��W�a\)�@����5�v¸:\���q}'����&9�ڐ�ut���6�FH���m�ز=������0�4X��*he�!:w�*u��ixэR!����������F ̿rj�)N�8�㍑ST�,k��a��>r����5����w���J
��Fo집�ǂ�Fߤ��ce'�[ƽuSfxL��'�C>�����mA��z7O0���K� Ǯ[N[C�Ou�GI��O��� ��gp�(1�tuu���?�YQ|:a�x	��|��lN�gcva�H�}=e����@YYY�sWi�R������+��������M�#���v�@�`D�Z(���".��eDR��RM"qFљ���.��̪��*���:��L�n3����#����]{l�[��W�x��+����;��A<�
�d+߫Z4�j�ꩴk��G���4L���qw�L}g]���c��
E9s�U��C!���'�,�����/��+�󘚚8zn�����H~���2�BfM\OW��/fP�~�f̌s�,�Hb��.?�)�`���`x,g3����j,��H��٢��E��ˤ�ǐ7N���;�����u�+=О��  ΃%P/�WN V"k+US��B_�S֗Q�{�K*�9Bc�����׎�r'?�0W �ǵ5$
�gr�_��v0�z�ZBc%�J�r��g�j�Q_9���#�����`+�ty$ڕ��vN&��/v �����S�6d�� 80��"�Oz��P�X���;��.|�����x��b}��n%�"���k"U*�Iy1&��2�0[#g��f+��������b�4��L+�F�ݭ0Q���.��q>`M����iF�J��{��I!�R��4��ݳ���31��J4`쉐W�k�c��pC7 )�E[g���J�5s��#���"�㔶�B�8��t4��\�=B�������]U��#�>�9��d�*���K��^��|p�p�n o��ID'�W��w�}Fr�#2���*݄,��Y����*M%R����\�Mh�6K5�ט��&|��Q��s�C��I�5�ū���MrM�L�Y!�t�M>�pc�g��	Z .��s=���^���v�O��ק�q�N�p��V)��O�z�����`���zPzjb� �NƸ g��om'�Ok��������h���}<&�T�=����"7�<k%�ۂ��a������R`�1S��!�k:������}�Ki��G��y��r�ouk*������g��,\2�p쪌�ښ3Ԟ<*Ο��V|}c��4@)g�j�p ,!X�O�xjLo�������g�I%����fL�0u��\�
M�u�L�ޑ��?;�5������VM1�D�G!YF�`9d��q�$�ɫ"F��k�cM`{x�X.��J����}�\a�J�z_����h�*�b"��e��T��u\�c��S�q(�������v:[c(Q�m���m�+�nk��^('���[��((�-v���e���_эr/�7��A~��Ԫ@����#C�AR�\[:<�rd���إ���E#�>2�P�ïm������pgfؼOe8d[�#�.�zB��B����sXh�2GϹ/4�'��]��l`�!����)�|1�y�܎��"��4o�@*��3��p��Ek��Gp�N�/7��6���C���[n��?S��� ���ɻ����9w�����@tƹf�n>v/eo��a"�8J}L~��d5./���X��TOؕ5�:;���������/��M�G��p!˴��q1���҆��a�k����9�����OVo,-��>ϗk��֓W�������g�h�i��E�8-W�S�S	���TE���<;*�A h���?�H�V9���H���M:B#:UJ	!�	Ӈ�pt�$�b������/���6+��]8�ñ܊��>ytI�A�S����hv���@�U��r7P��5�
�УZ�c�BѼ���r��������,���7�f�*r��-�������`�=�T��{������'��.�YP�i"CY�Y����+G*�3�}'@Z4�dR��$rL4�^|�3)��u,+�R�փ@p���,�3�9�a%:v��bO߶�vN����i�c���ȼ��[;����+�"���y2+�71��d=Bm�?\��v��v�~��r�3��̈́��Y-����:H�l/��[{�:˪�Cg��@Rt�~�Mp�惙�\_'�f!�f$��C�IA��i���E�i~�+Hfd�7ft�B��:��=���ކq��P��J%�D��!祎�\�~��F�\���@���x.��ذ�]���o�7/,�3�xu�bFձ?����N����*�(�հ��0��:T˟A5�S1�OMW�wPծ��=:s!��v�P;kʁ������!Q�8Vo�(�x�d�C�X���\XX칋�	ӟ���f���){SeiJ�Y���oȞǠt�� -��Lj��O7JS8M+0�p�~��]��t>e�Q6�0Ԙ[��|�I	� �:��C/��.�Q*u��ϵ|w��#�n�������+���u���� �J��~=�\Y���M睨���lǼ�v�6���g�ܥR-���vR�k�PI��]L�|K�=�`�e|�$�'�������H�����Ut��v@���?K���.�K���J�~-jP;�ݪP���<����,Y;u�ݧ�T��	!��	�%u|	jױ�]6Y�`:��P;:���AI%��%
�����ub-)X��{4�Ïeu����^+x*����2B@Cn���İ��n�D��D�*�� �Z���B��7�[=��������uS�Γ�$�6�#���T|��O���A��V�?��֩�.�#�6�������o3-�Fmf��άt�"e�z��+|q
J}����,����I%���?(cPu$y���z���>Ք9N�vW^i�b���B���jx�3�����ڱ���f�M��iIA�Z����o����-�Zd��ǭ��s�y��Ǝ��awf�m�?��m߇{)#�%��G~�K�1�&�/��}����}���$�Zr���μ���uB�����KJ���������%�jgtt�����\�N�@ъ���=�Վk���!7*F�,�L�K9�^W�F����dj-�#%�l�M}��֝TrJ�)t'A��R�..�S�7$\�S��vr���֤̯��Jw-N��t�:!��W_f�c��#���1ڮ�>�ü]�>N�9ڮu�e�rֺ�9ǅ���f~ܕ�$]u���v�b1��pd���+���9�rI��V-�)����O���sQ�gL3��nIyvb��U��3v�*�J
1
�*4%`�*+�,�<���h�w�q��=m�S8���atK��,UZ.����c�?3�!��;9���噦��vۚ�9����,��_	N���|F%��|9�.}1ƹW�H���&�t�+��b�����Y�&��MQڷ�u.5F4aE�N�\������֖$��Wo�l�,E|)Z[wU��b� cl�_ϫ�~ @�S�g�()�8H�h��gs�w�iC�x��m�ƶhk(���E����~������bۓx�o�=��z�c�Qͯ��=�X�zY?���_�U� �N�V�l�h'ͷ�j
������U�ۮ[82==�E���h���~�Q�[4���pM�
KL'��(M��=�%K܌����ivm�z0��0�Ж��q<�ݣ��~���W��{��d�_	�h��5��o�ភr<�CZ�:�V��+�c��L4��L�J䏖�7%T�1�{���k��S����*&QSc�Bn���<����(�?R��.���8�QJ��q/�^�<�,U �� L������Pf��j��C�b�-�^C��1���c%G���D�/�������@�����f�Z��,��*�9K�N��cӖ/[G�9�yt�	9�y��U:ctX�b�"D�"�옥�����85-�Q5z�ݤ畲ϤV���v�+��7�.�2Dyhkq���!Ǯ�C�a���Y��t�`#z�rM/����$)2:��[�O��O����n�a[D4N��,�p�3��ӧʢ�2y��͔xi�T�+����ГQ����8�y_�q����w$b�%�\�q'*:�p���w��OQ�̈߶-�AA�X�α2������/����SYB���<�����~_�+������i��AW��eI����;��A�,����	\��DBI�}~���x�_��kA��BL���D�xc,�������1�f��vVay����S�!fq�-��"��R����d�m�G\6]|��;⿅��搊��O���~�×������y��AE���'�M{s�ڃ���YE����.�%5Ǖ�^�V��4D��f䘦ޔ6���ڪԳg�������1i2���;*�G,�"�s.�XE���u1�՞n�n��-O˟�J:�x.w�T���5
���޽[���}��)a�a��o�i@��-ьǕ毾r���&�6/��U;G�;g:��I4¯wb�//�20������bf��C*_�hɬT��Qb�L�ad>[�mK/��W�"�mO�������3�������,d8�i�mo�>#�o�?}�f澭��{5o�����U����I\�϶|�`��5�3Q��F�T<�?D��ǿ�K��CH�*����ݚ??d�>�R�V"�6�2���@�Yk�q:����l�v�z�<�`���m��_��&F|9yK�G�=z��J���ѣY�;�f�D �anS�*Ź��rg��)�������9^QF�}	f���0!A�4\-09:OOڐ&GS�gSn9B��%�̝P�H�u��ɡfR�{�T�G�/�q�a�jg�mz�M���/>j�o4&�y�y8?�㪇.�2ݠ��F�������O�L\�v���膃�g��8L[f������	2��ߎ�l_Ҝ�p �yQ�C�{�CVE.CM�E^,On��h?\��p�H@���VS����\4�!v��6�A�զ,<FPr'B��!-�h�l�����؄	�qJB�,#�8�7P��L����6�怒������<4!�;���A�M۔�"�0D�6��l}g5��H�}����	��Jӆ:it[�K^��=Օ����?��ۮa�t���W�u�3\]�y�l�g�?�9�������4�B�혡\q���M
����u��gn&�|@4���c�?ÚZ��Q8��5�� �(
Xh""-`�� �t�	�{�P�n��( %�4��KhJ�KE-!�P�,�o�����r����}�/!Yk�yf�瞕�� ]>�������G�k�����ٮW��8g�o��o�u( �������D���ƾ����Do������ml�rN?���t�Yy�c�Vw���0��e�����O�	Z��ZW���'�B%oķ�'H.Vo�o�dW=�|�=�9��TPR�A�{�_m�'��D�Ir�m.li�ξ��9������%.	K��7�>[��a��[Ch�Z�m��#�K�<���J�����&�3�Y�=s+�G���k۝K|]���/4�o���N��E�ym��?�C�D?B~SR繶����&�J��Զ�e��փ544�F7+	r��� �����G|��U���K~������
��Y�5w��^{WW׿N���#��r��%a�2R�[)<t�
Ch��h�F���)��%��Pd��ERƛ�{�D`��4;j��'���X�q�SZ�MZ��g�������Y�fm����Z餹g���?챛��g[u�d6�6S����D"VW#�xc���CCCJ�NXH�㋖?#~!�U����[�
Us��n����E��х��[�s[�:�{�1>�7F��a�kK���]��[?����|�Gq���:���1�S�k��4�v���My>���2�{>kt-��]���S�H_��������u\v���38"p�O��V�4�0��?�6�9Ԩ����F���c�,uG;�wܷ����[���<�1�dLj)�׮�L-'w;z:FM�o'�<ő�?�j�?P���n�$�lvß8]����D���/ے�ʭ�V�}��L��=��tn��_���q�n�]+�q틸Y1��$n�ŝ`�M^�Y�u[!�F��4��|��y�	��\�)��l�ժ�Μz5��q.R��}_�?b���%⽂'�-..� �cpZ�o-�S�t���r���K�W~��׻ۊD�缙}Vk8�{�řQC�3ٻ}��YVh��	 o걒;ϴ�?�i��57�YK�J��h�[���Բ\wH^��*G4�P �����!���_�ۣ~���ߔD��ZY��o��
�����P��sQ8���Y��9�/��&�L��.xݍ���� z_Ǯ�ō*�^ �s��wO��P���}�<i���ߚbD�6(kg���:᯿��]�J���i���h��m�K�m�n �e�X�&	�g��[�.>� �ڿ?@�k����I���5�-�!�3^�oEW�E��W`�$�����q�|=6��֚��F^��]�A�WU�fDHz��Z\�(�N�
�Ͻ�9�E=
A����Ӣo�Z�E�,�>]���}���E����ls�TL�*5y!k"gࠎ�U�70����C�q�~u{�S,��h������ڍp����f�E�(�n;,D�7�w{A�inE����n����Bz����(�s3�x{�+4皝��w�5/X1��ٴ;�������#����W��k"9��^@8���}��5�`+T���SD����

��SȨv��8��g�l�J��Z�(ba��%vW������t���;��p?�(���e�^�CKX5{��8ב��CV7�(�v���:Ғ7���zS+�0y�o�S���s�E�dI6�,Z ��g(P�V��P����E��"O!>(0w�ϙ�΅����������-6�w��L���n�9v�O{����m9wo��ۉ���߿�K���'�.�g�?#����F�3����g�?#��F��3�P�y����ċ�'�ط�R�6��Ijut~H���	����4M�XKN+�A�U� ����i�$a�d��I���"q�諩�7^��z�:��`��m�J{��^^a�;���R���53o��8��Z��Q�2�%���I`}n�/��ל�[��*����_����{��6�}2I~ڕ�V���oa�J���H�~�_N>�)�^�ql���������O�Jb�_�NR=Y<��Ю��k&�p ������ژ����.�pv�Q�7Y���T�&Kh�Bͷͣ�����\nU8��T�ʘ���gB�.5�V�����W��j�˯GJ�r�G����������9ݹ�V3��C��ek��7����멒ٙ�D��j�P7�V�tO��&E!CJ�@���9UW����;(3y��1�\+���c ���V3<�s�b����/-+{��kT���P�J����gB���	��y�颡�7ɐ�t�
=���l�S(aSA�Z3��mfK�o\t��Q�P�c�wU(˞�y�k��FŝC��`"ݷV�d��r�:�:�F9�*]�� T=��'i�R�j�'Z����#ز^p�
�->'�#���)��se�~���g�.r�`�w��8\+�\��������b��4�:m&<U��j���O���f�\��;����{_D*rO�c+�ttu�D;-N,��`�����D�&���&��A5t�x"�����_P��aߓN�/��O�9��7�{`��I^��R�C�^�c�W�
i|vltAS�;|�����򲺑����A��y�?�3��knetyY�G^P�a�*�<�Ȅ�E�H�q�8{��b����s���e��K�rǟ�e�����p�*�҅j������SoX\k��d��ܔgG�M��c?JB��s��<����t%w}��#���v�eC���}��i���$C{�N�5ֆ������}{�L�i�b3n>�`�!�a����1A�'Mb0..<���Bݽ?���c9�����D�K#Z�w���$Sg�o���� �rhd}]Se�k�R����<=�:-:�ޣ��3@�zT�	��k�SRo�����߯�ӽ���f�%�T����ȸB-7�$�c��aӒRR�0���2�Ҕ7J_/s�\۹�0dTIT���t�c�K�f�f��]�d�)��7��K�V������X�pr�����nX�k�K��juצ��&���<r�d۴1�����9���Q�|�ԑ�Y��d�=��E4��lջ1c*XgȨ���K���Cy^E|�r0��k�a���:�P�7|r�f�ᑁ[��N�TUi�DOEjϵ�;�D_ǜh��#�Q��7�i�l�TŐe!R�9��R���<��.��V���-�e,֙X��:,�g��(�wؖ�(�ԫ,��\�RxP�8�3���'ɞ�z9�9z���TQ�P���k��. 0u����P��Z�u��j<5m��P�?�$��6s�7�H���q���My��	��Í�m0�k��>:���o���
}]]vW<��}� P<==�Ե����'Ά]�pJ���H���'�{g�U��@+iʃd�ͺ@d�NC4�~A����G\�VT���`|JM��~1�Y�-ڌt�����45D�o�F2k��-))��g�Eo�=�n����>���A^��t��6ǰ ����K�_�m=�R]E籢l��/ь�<��EIE��xui0:p�&�Z�E]���)��f�;8��H��� 5%��5��NI��{��f8��kv�N�H.��(�� �q{{�B�����L'ozKW�f� �P�D�Pg9��
j��&�����]j�~�����uN�B����W�Z�x�����9�h�Na���9V����^�.0�Kqi���Z�����]�}ֿ%oF�ɯfXv�Q��� �X���|Î�К�0�]I�	=��h�M!9=���Y[{�I�������N�n�@����|��y�^h+��^�@���V���,�rWY�Y�%�ע�C�F�ã�
��P(Z�@����W��{/@�AC�">��I��$�>'a1��qnn����E�=�<MZ�T�P>c� HN~ ��%B�6����	�2���u�ΌP|�5���l���Jo�؟�J�`�4��R�qr���B�k�����P�VK>]�r1]�q,��������	oUE���LH_����h�~U���`%<���j������'�ʿ?]�G�ru��:,t�a����J�Gǡ�O�����DI'��⌑v��y
r����п�y
T
}�<d涹�\�E[�gh�U���2ۧ���Y3&�X?ܜ�#dh�'}怉�D��I����xG7��U#L�����5����x����-aqǰ���:p��5 ���eޓd�3c(��5���`hnd29��\*'&x��e?��t�4�-�	�j u���&!B�����H�8AQ�����_i����Ʀw���X���ZC t���9��>4j�@���oo_��w��treH @�P�������
�	�b�vV�B���n9g%�t��G^"���oD4r�����q�	�QFX�3Wo��R������ߍS��\�.��wb�GC ��)Oi�6���m��cSR��|/uo�D��r���|�@ h7td���ʆ@�����G�{�!�jTݏxE���P䌋����|4�0�uLrh�&�c�El��6$Khh(�������Ƅ`���n`�9���Ŗ��ݧ����wϭ<�9eS���ܬ�s|o|
N���(��U�%a�E;�: ���h�^R�=X���W�&k�U��酼o�������
�E������?0�zI��p�^0(�%�5���䐹o�)�����������6�0�|���Q
��Í֩�	(�g�>]�>Ud[�o��_$�!�2QGC>g�)~�L��k�@:�.;!�l��a���;��j��xM��~w��̸�Ǐ��	+˔~����d�s��D�I~��CO��ϸ��f���g,l-��I��u+$$0eߑ�AX�;KO�bn��� �	��^��CqY � ��/m4y���/H�������mr[0�_��aq�ܙ�A_�F�Eg���S���G��G�y?�л�,B�:���#`CLp"����gUg�G�}qk``@s��7�i�!��`�/��ܙ���NO���t��#��mG�B�@� ��q�ٹ����[���~K���5{h����(�^3�}�7N�����>��ty��p-�L"������d:{J�:k�6�������:��7l�ۅf��.����~B2V-d�/�S�Y/f\�Hp�D�SR�12޸q�0�+ҹ��,o��r�g�5�/H��j�`C�Y�Щ4���#����a��7�wtlݽ�:B�;�j%�$��D��*R�x<M��%��Z�4��"%�~��g5W�)]V��=-J�S��dP�E#1�PQx)��t�Oޮ�`��#�0lE�z9��i�t/�C�.��&���aP*N��=(�޸wu�;LP&�m,f��~���ZT���p!���~.�-��{fv�@��u&i����O7h0褠����� ��A���E�v�(��[_��L�"ѓ��������FA��H8�i`���F�sc�3F�B{�H$:NX�H}TD�+���C �0�	�'F����@q�]���v��u��Ӣ,��ŦbPdy�9Z)�mn���m�x�����n�S�En���������g�@D��ΠZj�DTb�)E��O�D,�<Q-� k!�C��""[0O_9φ�Z�'�o�<7`�A���r��W���ߊ��M�c��
� m�����η~�f�"�#�����Q�$��ܜ0Yt���� �$m�mI��"Q��j��%m
��zbjd�� wa���4�8J;�Y����%��`{�h���X� �hP	Pq��8��ϼaeD>vx{��J�1��>��ق��~�*�AܕsV</a��PZI!\�5$�����Ċ�ZN�\T)��~����ip���qg}����Ǧ�b��"ш�1�<�P�|<���/�[�X���W^�$m�`�2��U�#�J��B��GEu;!R"8�yLƫ��8�ķ�&)���4U|Aa�:�ͩkc���kX�#"����ƢG /�Տ�i&/�K	��ꂼ�|i-++�x6 ����t�*���	�5���JR�1�DY�v�F?+BJx+�m��w���S��e��<���'�A��N�*R��,��W�����+�Z�h��Q6� ��x-940C*��7�2��3v������;�RC�a�q`�j�@��r�f��xB:�wӻxX�R�	$[r� �B�(��`��~� :\.�et�{Z,\>�|� ���/���� ���UK�V3G@L�ڰ�p�6�������Y]�:Z;ȍ����{9F�B���~������XlzŶ��uv��W�ώ���=��U���c��������J��L�.0��f�#���~��j�j��v����3��+軗	�rߤ�_Z��6+����Z��d�Q}
�0Kx��Vn?���^�o	�M�0�#�Tw���:����s��x`lG�(������f
<�z)����6��csCW<V�4FZ�ۛ�;�+
�J�� �͸��k	)`���j�O����d��?i�CW?�f���d�d�� �Rg�h:ҥ���@��h���%2�+GAL�/��L��U(Ƶc�$�eZ�K�$�t���s���b��pl�Ed~�ǫB��y�I����XVT0WʁZZZR�����P)K�;�\<��&�QR&���Uj��/���th=�ܡe%R�@2���Vd[��h(��K�u8��\�J/Z�1��L��U _35pXC����l�0�4Bb�z�MN����hM�<��)�\6<��0����Z���i[A�*R������M�1�X�m�Ԕ�E�#aV\�ΠrS��4̥��Ol��z{g;k��t�F<$7u���{[u��@t���}�j���nA<q�5��)����EG.�Z\�<�(Z8���o)��fvܝ߁n�sn�.|&���t���\1�s?�=K���bW9U~��4gi��'5G��b���3��C�HO��Ԑ�B�!tO¯�6� �9�����γ��Whm�T�SE��τO�\������cc��K6�w �� |�д��q�D��Dd���
�Ʉ%;�Lkޡ�-1�>9�Q����x�y$"��C(�H��$�Z�,��	~�P9����p����:z���!A{nJ@5��ڈ��8oYu�E�i�u�;{�aڙ8	�����-���8Ø�s? �I���CE�-���øv=�b��OY��JD(=9ɹ8칂z7���q8�����Kx�f?����
��EW�n��s���t���t:��A�;��>�)N���N9�":��\�󙌼THq��F�K ��?<.B�>����tR�!{
��Ru��4:���8z'?X�~��Q>ц=[�J��{��9�A�n�ä^��X�k��5�ǟ�1��i�*���u�aj�7��ɨ2�҃te���v�y�L%5'����e�������,y�twPO�����w��;��?K�+;��l66<��t�uw�2K���Wx��k����:wS��
�����:��.��&5c�o��9����1�=���u��KT�̘��i��f�f-��ET���ݢ8}p�BݕE���70m�Ag]�O�0�2�gs�ƢSw>UؔxB�욦�����j4��J,�1��v��XhݬK����XqO��|�q]�nY�@Bt��������h*0Pj����~ց����
�UUs�cߜ���<gϞc�5�Nv����."��8O6��|��E��K��#S��a��}d���� �P�@�P��xL�����ɜ1��򏎿5�ml`,�92���L+b$87�bNώ���u��n���I����Y��$~�F�+Is�H,���M�zGv�N���M���O}&�" �	S��W�?�x�͞�����Y_X�>�$I��q�;Ch����,O����-���M��K7��������={�¹|�b�wQ����SB�<z�-Y���grk�8�mx;�IB�zO�4}�q��!�2�tl��eS��B�	�zLSb�cPu:��R�j'��b=�Dy��꼫��DON�v�\,��Y�iK���K�����_���@_s���~�J���G
��ز���D��Y��&to=&U3�{�1����	@�<� ��N��{�=�l�a7
w�$�3O�����t�u�y��߻0My�6@M$vOs�o�Z�JZgsnME���{/.��z� fR���0jV?����������c��C&�Sɍ�Mw���>�`��o�P�J�}��Ζ*�Ň�%�����N�V�!�(r#�s-�u,��/!�MR7���h�8:w�V� lhh ���[ �,��>d��.�\�A�,e����d(��%e�����Ч�Xy;:&�e����~��������G�f�vϧ��N�^R<���`X(ђwK&_q��һ�\�x�;����`�x
;��on�<���D�d�HL�k�;��41�(�[YBH76v3�ӱ��M2�M��s��UD#�T�T]�=]�$�e���m%�A�	<��W�{�:���Z��Nv��˟�G
����j+�?�������_�>�t��By>+�7�bz��X���{"zȯ&,���K�?�Nr�d����$�lQj��G��:>�5���}�ΔXZ�\bXh�~�p7���6�8���xa�6j��B��y�˥�1ձ�c�F����V�T�����R�.M��3�z�7zsq��ۥ��yv��2_tu�N(��^(��ޔ��q?��\��/�OjHh�7���l��5yFj{��h�@X����p������}�]��g�kYj/�����~��^�{4j(�ٱ��J�A�,��A<{�x,��W ]�/��������T���k%�vQޑ��9����E���R+.���u?C�̭ŮФ��r���`�z%q����p,��C �X;�0*%�������D�K;n�����J�C���jL��^�|j���U��L�ΑM�q.x�!#�'����b�3���.��*H�~�1����l'Zߨi�xbx��}<�o{9H;�Wr�*��2\u�|��e��0'��Nٜn�y��x��w��ٸk�0rZ���т/S��ej[ZB��>�gp	)�`�ˤ��ӱD��׳���`F�(�<�"I�_}'�?@��2Z��������/�Z��w2��\m����b�S�;o�Ƹ������%�P�R��6�"gړ{��*����/�_�?��^�sC�̽H�����cB,�[���ޏ����R��Q��A��8�:kp���8D�+���]������S�Sb�)z9s�.�>���C?����uI��-�N8����]ɳyK�͞�� ����=6;�^7)�����Q%�AG�x��I��)��U�+�(l����SY�W.��|'������%�վ[�;��ݤ��cѢ0�x(V��5X�c�榀Q���ǣƙ��îlMQ����&��xO��h���̈�(�#�Æ沼�=\�g�U2��^�a�(�Rk 诗���*�dف�'�ܳ�����X突3����}s��U̐��MoPVf��F�{�W���f�%�f��d��{fΔ�S>wZ��j�w@��X�ܱ�7�Zd�_{��Y(��RV,�?��2C�r�%x�-{	d��	}�Q/�����F�-Ϯ��ZL�^�'.���qq�T�T��H��V���TO�Қ��#���������cZ�N��aѓ�]ސ�ja��x&�Hn�=(s��}Rm����!t��_�>^�����% �4�b�!�}�N��V���_�
�jM�R��Po�������D7k�` E�{f�����dzJq��|���?֒�j��`��rn�cr���p%���W�I�6��+��7�����<�y(r����ڦL���'���T��e�{h/=���5Ra��9ob.����*{L}xDȲa��A`�Q��Qq���}8�������W�(���o%r�`}Mf�`ݻuA[5��l��\B!��p����8�L����c�l�/{ْ��J�c�":���z����!���2ǵ�w%s+Lb��ar�����g��w���Mc�&��^L�lP��j�B6[\���lQp1�D��\��u���V/�Qz���%$��IR<��v���/������a��a��F��Mqa��i_<~��0s������Jؐ=����_��&�:��p��?���� ��/�����A뉟QIz�J-�/L�����U��u��^�[~/HW�$%}gn�x��}���=��� B��ݩ�/^��G_K*Ny��o���.��>�����L_����	zh�Nx�L}ޏX����9�
�xʹ�a���
a���`,讅�N�� E��o��c�y�4���hr�;,��0��z�O���6̍DV��H\�أ����/l�����P�y x���~M⫖���0C}j�� tR�T��N���Ř@WZ�[N�ck�!���o�Ի���κZ�g��0C�荎	�����i����f�ә�Th��©A�����<�/���e���;� Iヤ�z���ز��"ts�͕0�P˻�E��`E/���aW�U���[\kQE�hш��3��
>FG+X=���v��f=��k	U�Y�c-w�=��f-�0�60�6�l%=��	b4���ߠPۧz��6=åƢ@�eDN#��4�6!��T��&�d7�;�⯌��W���.������x��54���4�y+X����8���Z��:\0lU���S�#�^*���n�����g��:�>*�D's����"��h�d2,kh���Z̑�()>������{4?*r�1��$����������_x������4]�"��Gzu"��Wm}���2��#r��<}�����s
���*}��kg��c<��&� ���c��������\�Q����$��ɓ'����1����t�z����^�������ɫ�O�N̠
�*�F���d@^@0�u��Q(�k��'D�������PnII�D�z1=��ɕ7��\Ԙ܈�g���ڮ�݄]�Bk\��7�9\�q#��������fi��Z�t��%2"Jd��4F�>����έX{��z�ѽV���.�>|�ނ����z	tr@Nfltt��7�_4^�>� {�P�-�qQc؋��m��˜��&9��J{Y�8��Tܵ�WY��Yy �u:�8��o&�� :(9�VOd�]%����J�����[%2�0�3�����l�
�ʓ�S���6����:��@�bZ��Z���wQ�ǐ���Esw��苆g��嗱�
�����
d��������?�#)�Fi]Ē�욧�NB��{�}��,�ћ7��]��y��2P�Ott�t�#&"���:� Вx�����) ����VK����j�G0q���6L�݄��gpP�s 3aQz>0ۤV� 5��{fX��y�WY��L~������	'�P|AAR�D���D���#�FFw	d$�f� Ul�\�X�R�����ojiy�}DD�m{���[lj�9�,
� Kdt����h�ĕޕ�w�z��y%w��JD�4pw$ƼkQX���!��%��,�5c�<��:��ŻC�.�d?�:�_���3��`O۬���TTT������&�8����̉�K�f�����C��@�
|y�&�2��o����O�.ԶpA5���idtF�[��66<-�A�Z�δ:����|�RU�7��^�k��,���D��B��B��Kj;�=�V
x\DӘj�	��%�	�"Xj_6�<��K������/�ײ�pts�笽:�I��K1˹�}58�\U^.�O�i�r20���U?;
�Q2���n����OI? ���=��4'��Ʋ��F���,g�ҿ��T��G���c&9H=��?4��{�؊3���t�l �[,MM�7��*6��;(���.�r�D�miQ�MN�Gh H[�͗���v��|u@�l�Nw'Z*Ox�����gkk�*$�
C>nt�����k��u��<~W�|�4��%OXӘ���Xa�"�O��[z�Mo}�)'HU��#{_h��k�h���x�����ʿ\]\䎽����q,�06���]���^��72f�*�0��20##��t��%{�]����!�f��Ճk��]��ߓ�p.U�|�{{{>�2�^�zR������b
t� �"��M���h�6��=�[Yy&Kݒ@j�(4����M����B7�����x��:|FN�Xq���J�B����?����allH9��9H$�7Fk�r��(.���9P)�C����G��h��Mc���� ,'dee}�3p+ ��?���P�eM��O���2;)�@g�`��ȏ:�(�;��E������5�^�����v+�
�ȵ�m/�N���dr;�^�F�b��g2c�B{e<�*"���� �����e�Kk�נ����0)z�9>�����E7N��W�
F_[�1�t�ׯ_�S`�_��3pBF�&QjA��e�_��J~�rA���|^g9��w�ڔ�ݛ�a�2p���y���ٟ{{}������qY�s���lgg���̕_�
��}x¨<�vD�����*	�w��ǩ�8�~u~8�7���K(�Ӿ����E+m����ZZ�;[�2�M,F��g��J�(Z�E�c���ň����t�=x���-���q��1����*�%8\?�{�7@=���$�"7S``�z�r��O��'����� s�zFp'�[��iV"����r��E�Ir�WE�"��
xP�N=}}��D$D(XZ|��@�Rjز���	G��Q����)�1�q��`>��84�V_�
+�u��m�E�R�R�2x�h� ��(o��a�t�%m��(�c\Gt�ʌr�v0�D�~?L�u�^ŰὭ����Ooa��`��-+W�Q�_x�2�<�O�^%xT��=.�~67����C3v �ƚ��ʧFQh��\,`x�r����a���f�K���j$n�� ��̬�`�%�o#7�L�Vjf�)�hM�e���������4a7W�3T����-�h���א����J#��b�׾=�����GEՌNQ��֞�(�Gh$@TA����d4}��ůI'Ckk�)����Y�#��4U�&5
#�����AT�s�vϊǶh��e�6SɃd�c����G&''�n����yj�m�(�1R&�Rq�P����E������l/�jl�"Y�y�F���3�"�1:�j�'��j�R��?j�,_��~L{}��@A*ݛ�a�%�OA��ܘ�H��i*�C[�bؕ�����l̡���nh]��	�N��zq'����"�&h3K�0����� j�Z��xJ��AJ�v�?���QX�Xj#�C$����JKK��4�p�?}R���aY� ��(�e��0���,�8,��:�b٢P��g��2�:N�����z���?rM��:u��3��P/�+J��5JJ����H��Q�2��Gqqq���9�8r��cx��%��iQ�ק�������鞆�F�z%�i�<�Qp�GQu�M�>���{�{��������"���r"��C*�'�p�x�g�N�;Uz�<����}�9�΁�m�In ���f���j�F$�-0nC��z��j<p!&󰆽ZF'��63��7}�0��
��S)=����n!Y��Z�s����
v�k��FXi���/��o-rәNq?s�@�I=�aGϷͭda�u���_� +Hu�������	w���0U:��:!z9��R-���W���Y�z/����z�7�"/�ZR�e�r�
L�=b�t�L�&�&5&��@��&t�$L��eq?�r��t���E�O@�f��_X�f��	��z�����Q�q�Q�L%�o���̀���z�\�T�����0y�*�B�������̚�L��}�9��N@FQq1��6�Y>�[Ww������{��k*�a�M1���^���t���&��-��v ��4�9A�^�9`ى�>�!8�l��h3��`=@:�an	�z@qD܃�Ku���(�>8���y�����8�Ǘ.>~~9HJE�M1�w����_����;mZ,ay�{�0rO��(%'�XM=�En`p��/+�v�$A�9|ۤS�w��H4Q�B��q�8�raL�&#�L���uĦŔ;0
����/�^�����QyB�!"���9��߇\xN��,?�M9��(�oȏ�VF�5ׇ�.|��)֡t�&^p�I~�� R�"e���pH����8˫r���������r������H���]i��7VpA�"�Ks�t������(�dV�I��|D��c*�*R(��F�6���,��P�Ȃa��I���g.>�s �R���k�"ѹ���;�v��{�����j������cSL��ʜf�\���%eێ���p���1�O��QD���*Z���%�\,�4�[�8٫󳪑7.���Z�2�C�t�V�
�)�!��j�1_��ȷy�N3�_��������LL��i���D#�R��b����i�]�#�6�"88 �	�b�<+Ao�	T�����؂�o�������>*��Rc����x���X<�(�0�uX�AQ���:�Nw@�вw=rUۈ��i
��H����V��>�\�~�RŔn1�X3�R��~�v?e��Xm�tl���i��	����/������SPDدQ6ŧatP"�'�4��x�!A�}�G	�;+&=�]Ƅ�y�\fn�}�U�C�I��Y�Y�0I=�X�*����nP������ �{��r���� �2s��Ѐz{s/]����UfM��Ԛ��0+�,���h�������`��:_F��
��> �����#���������iR����'����=є��B�LB]����%�g��ć���3Y%�
zlA����j�㏠shgM�Iq��c`~U����[�(d���W~����^@O~*�$��U�c�\�� ���!Z��ܗ��#/��K}��a�ϝ@��84��aL�ҡ֦^��"���Τ?�R۱�(���9�|Ku�@]Q�zy��ep��7�
9Hua��<����
�WɏJKŨ��T(��0�� '�:��
�Q��;�:�P���i�Ն���c(��o�Z�*3�T6�{a����$/���&���}���S�V�B$é�� ���.`p�yЈi�K,����IA����}^�pcek�t��Ɇ�4��E�@6�.@���� Ef��+82��rw|\P�/��Q���,3�hy�Q��'�˓�%87�}\O"�Z���]U�/��38�f�B�V�H��ϮK�$��[��)��qd�\͠�i�.y�V}*��=�(. O(J,4��У@��`�I�W�T�d����N�l׻��;1� ����Yy�v�S:H���bD�ѣ^`�=I��i���c�=((�E.�3�_�T�avB5��r#��H����ɎyH���v��_g��mQ_|`ݞ���8�5�q��s�msk�oH�xh/}q��[( �O-���Ϣ��By��޻�����8�Ȓ}@�y���j���w�"�7�������ܿ�}Ӝ�.�%xJU��<2���r���|����N�ow~��nOX" �7�=�����������|+���6����/!q��~��S+���H3��	��w7��j����>�JlVMS��8��}��6Ҋ�Z�m�^�Z�m�W�r<��A}�AN'���3� T4)~�NKPyRx�ǧ;8Mm�$t���#�ꫡ5a��
��{u-Yy�y%�:��8:T�Q+a�)���c�<�\���-����࿏6���8tпO?�������f<������g���f�����=����e�W� S)Y���-��l����������%�b�IA��,�G� n0`��Zٓ�	�O�ޠ��F���T�Ce�a$K�%�^������oM�?��z�Y�;��Ow�ٜ:��D�g��˟<_�P��}z(�p٦�t){�ѓ6�Õ�i��>�j����8���٨uZ��+���;����Nμ��-���o>q�����?����u�#���T������[y�N��3�X�*R�c0C�&�y��tp��	�S�}K5c�ZΥLt�3��~1as�g�4Mڦ�.�X�d�$71':=������z�#����:���B����arO V6%b�ڰ�ӿ=f��1'�&d���.�Vt�乣�%/�B�e�b�Jg�Ts����J(C�ǳ(Aul�RǬgQՂ[����[\;Ժ~��N܋֌�ĭօ��N�#��`�ׇ�G�v?u}�V�~����m��_�3�Xd:�x^�! ��f���ٯۈ|���\��i�������'c�LY�ڼ%�������t��(�co��1s�i{or �s՛���\���\ǹܞ��Ѷ���C������5�m�n��������y;��[�%�wy�g~\������1�:[�}ϯ�C�
���}W�m�d]K�r�r7G`�-[ �#T�5��r��+�T�+�$��o���E�������u�
!��3gX�����8��]ժ�`
�L`�Ė�H�R��ǋ'�oȺ����8���4�w��m*�R�RG��%89/t��40<�z�3�%f���2!��m��mH6�YN5����8��'��EC���#�ċ���.��֒�|�r����@[�Ê��#�?[�1]�+3}f�E{�X.��R*³5����
��W:�u_�3�|ТŎ�o��]&�_���}x�%ޑ����"j��G'���Nh���q�W@@z�JDS����{\��Ű���枞Q���5_���P̲&�ͺ*ʲ��W6N�����3���ɗ���;�d�[�%�T��-a�2n��0���ЯCK� ��Q���:⽃�.�f�i�]��f9��>m�)r߲�K����ҝ(Z?\�gdl<vj.?����qΈ���5�A皉D�Vg��4��c��=^XmH�bE���"ThX6��K������߮ﴟh�	|�w��u���#������D��||�k�	�z��5�{ks
��;q�Z�d�M�;J�{r5B%�|��-j3��놠&G�Qj~
7{�>v��d�H���-�%�x��gs!��-F��n����ő�����*���??D~���8���N����$���^��\!q�,=�� ����}D�Ć%R�'luO��!W=|�ԕ�e�iK�	mO�R�����N7t!�5=�O_ę{�Ǒ���뜻u�w<�����]��K�Dee�$r�K�w�s�G$�oJ.�21S�_�8�,����;�&,dt��x�N��-q���~d���s++N,H��N&�%\O1���3\m��X�n���3��D=�Wc�w��gAn��ۿ�s��r�^άyJ�~c��1�rc�ͨ|BV����r����ɺ�i�H�<G0m/0[I�-!�<F�I&Nx�fo\s�7��-?溄�)�K��}��4\�r��t4A��W�V?���H�	l�� A���m��)�3��
�6e�)%��G���u|6�����g2)J��mtZ; a�_!�"]V�:/;K5������m���An)��&21��>��Z촃{���pQ�"S��{��������Mj�HZ�����������Q�A��PPRB�i)�J����z�nIi��Q:���c���眽?�}]x)�g��b�uϲ�]��9�Y��$���v���1����7P�_���`���F7c	+�F���ʾk>���V���"��t�/y�-!�[˹�K�ġ���D�Б��cU�t�V�l�Cz}Sl��1��2��;o�"�p�|����7��{�Z�<֢乯�n��[��Ю�f0����tTğܸ���Q�5D�i�U@�\N(w��;h�
���0�@!��1�~a�B�8ϗp���B%�ت�5<M��5���]��h�D�(Z�`�Ax��P��zck��g��Ci�G�ই��Q �:���?�&�䓶<!�P�����Vb�F!�����x667W'ˠ�ȾH������7��X�ma�^-�#zP����2�Z�lޓ��lbMA�!n�oi#{3����f��6k�D?��_f	`}%�c	L��~sr�lx=P�F���NJ��u|��?�{�W��3���VҽfN-����=;CW*3��^���a+yw�:�\��̹��i��H���6>�!�6Èچ죛��e��M+�7�\�\D��V#DWb2�f>7�����C�#��~؁��p����(�.����SlF�
'F�`^������v�Y�3G�:��m�^��S����Ϩa�y}�0����Lk����k;�`�I����{��&%A��An���:w��^�c6&�\�"(���l֜�|w�l�����!�B<MRP�/�DK<nZa��vx6j�"�������,���v�t�J޹?��۽����@����2b�ҽ[����s1���'s?�+��5d��P�+�Wp�)8J���<�;�����e��xE~����@�&&�M>��B�:l,FU���v�w��}��M>�pd-�����.3#��ejb\�H��Yo/�RY��`�M��t�+��8\u�7h:�+�sh�r�_�1���-��e��j[����A.iB�q`�
}�X��f=Q���Lm���S�p�?���du��/�/:%���-q;�:��ݞM�lV`��T�]�k��Ih��®!�k<e��̷�t��U�[ڸ�È��9�a\�u�#A�݄Z�v	ͧu=A�Z=w~���$�i�H��@* �ӯ:/�~��O���!�?a���w-����69�u��J;>�0�8)�u����Vϟ��(I@o��8S����Ч�&�������3;%��q��^}0φ��f��]�$T��{�o���9/jj��k�())D���_��0� d���۫��p�1�kep�a�D�qZu3�G��и��h3oiE�~_���a�N��
E��������?�[����"q�N҃-�Ӄ����u��:��L��z�s��]U�6�>`�-�@7j:���w
��{>��C9��IHZ�h>�N~I�>�)���ֹ����{dx��*)�:��4A�=�l��"r�4����O��w^��i^)����h�{{�#$Z(�!�5qIkE݉���(.X�����#�*�H�]�堙�hҦi�\ۊ��2(�c��-�<�<�m��GE��҄;c�OBׅo��{�A�c�F���|����E�h'�ɬ�H�5ٙ���_&�)B�Q��j!]Kb��н^('��
��}��& z��o�v�Y�c����R#�ת�̨��F��Bd��{������g����w+�}��*�4���+�b楏��A������*��*�n�f��DRX�Û7oV@�|%�����R./�Vk�v5�=w�
��e�3����^F!"O+��ج�����yN �z���#}��ÓvZ�I�n'�<��T����z �:�Co�r�
R�mD˩&0���IH~��S�����Oޠ6w�re�E��x�D�q����^Z���h�u�8 �Q��[�B'l��F�$(�K����OS#��DV���b�#��!��c��<#|��%�g�c��/wL����(��u]B��q+��_5��Et���t;�,Qz3���t�غ�w��:��ֈ)�K_N2w�I�j�o�)qCg�u�2"�,[m� ���'�7�`��:{53���a��Wm�������f{�҈Av<�i�4	�b��mippG�� �[AF��\���jI��y� ����.��&4�(��ݨ�n�@>8��}��)z��p\���#�k�r������0�Ƴ�-�J�{蘙���m³ȱ˕���$+q�����[�2�i��]�ZO��-l��­���0��wKzԡv���D�����4m��D��V�]�w���)�?Ox����H��y�AY�B�n�#��Ɣ�SJ\O�5������;�������c��c�/�D��(�������8�/�=�c����8&�F̭bn«$^�����͕<f��;N[����I����������{{��dA_I��Г���Zb�=�ݐ-����K�U&G�A��%� ~�D\m�/��,����_��߱���<f�_*جK��~��VR��y	�.B^���&i&v��#W���#N�9ی��MlX��g�13��'��ʬmYxm�yIT��ʢ�a��eǴ�����q�8�~�sLݑ?���B��6~��d^\��;�>D�L�����Kq��@�#"��=溴�����w��:��na�X���)�]+��z�a�j:��]��Q���L��-�%s<�j�a[̓?.>��ò�_i�ѫ����FP��+�+Mn���"��l:�"@���H��q�su��JKBQ3�Ej�A"��OՄc�C�ĝNs���P�,��0	����������lbĠ��0A�V�T7 %�M�%�pK�]��2��z%��!.���������|�g܎��i[��R�~�u�gU>D8y[�C塗WS $�%X+[ѻ� zݮ��(}��s0����Vt�ʡ���q|Y=��������Ev���Ν�#��mF�Wq�� ��quM�M��t{���>V�y̻�ٳ������o��E_Eb����W�ם��0d�ꔒC���i��xeT',�J+��_U>fI���T�����c��%koE��o�aj�-%_q1�8�+�>�f�j�Z��V���0�z�7�sAB�� {���޸��q�ֵ�>�CE��E���o0a,ikɌh`���U�m�3���V�'�M8Z��6�_렏�Г�?Z//��*j�:�z�������i�Ԣ��Q� *��H��|]\'5���#z61����C����	��K����5�¡Ew�y�����Ԋ����=��]��։��e��7a����=��;�7����|��=6E��'��f��ry����Q������1zo��/��a���9���4	(S�ZοJ�K��_�2rom���*|S����?_\�'�{����"Ӵ��'{!P#���h��8W�G�k�r�zMe�>{�_�!���XZ%����.vb%�mb�e�����K�-��,zuJ��+����a�E�jڡ�%�����d����a���%�P�ŨaY7�wdߋVB�F��N��q����+�� ������mѴJXNu�#�U"��tӎf��>������`7V�yq\v��\����'��3sֲ/a���bx�D�A~���Fv��~��Qat$����ɓ8t��p�<�k~e��߯V���;����%�B)��^s=YE^��&���Q\�����9�A�,1R[�{o�l�0|��gK{�����ی�g�T���_`7�sssu��~�*k���1����<�6��9��2=�C����>����f�!�R=es�������2��-�����ׄ�\����������D�=���)���Y���N��Oג�~�����2����9�9�(+.�B�!�V�=Ά[�'m�X2�n� �ռ�EI2,;�Ƿup,z��F��H�*�����ltgR__Oi��ڷy�=�>c�vٚ�ڳ�n�c3uQ�[���^�]Y�����X ���Z��������-��e�bc_t�����k����a�yX(G��XOUhw���/��ǫ��Lu�U��b7�������U.˟֞�}�]a�.�I�7�🟬��p�8��Ǜ�X:�}a"p�e;(v�naj��t�"��w�kH8�pq�?��������krrK��$?X��=�8���6
7f�Q�Z3���
��0A����'�J��ݝZ�U��=倪X�<~��Q!��.���v�j(�H��m��.���߿)ݼWz�?ji&'ӄ����_�����|TW�/�D�8:�]��
8sMȗr�_�'��Z����¼��j[A�p��N����6�D�k��>C$>�mBG����Zr"�^�}�����i���4M̀��+	���Vq==��{߶0�P��������ү߿!��S�ȼ*�\%|�����|����	=c1p_p�ND&�56>�c��}<?oP�[u||��]nbѲ�R9uu
�����,~v��@.��N�������O>/}���N���|�A�_c��Jo�&6A���Ȩʂ(�0 ��DST���&)�/����`z9yy��tX�T4���o`�����/8��Dh�A�nB��cՏÖ����x���*\���B�>!5HR[SC�{j�/�4�k����M������E	BDJ�?�-t̶���@#�mi�=mi짯���4�G
Khw5b��2Yr`��\�JH�^K_�� �P�+z�����ǭ��efe1Y�Y4��A�=,���?���t����9�M��	�t\	�"b��>��ro���a~1��W�on��*keU((.�QS#
Z�]g ���T�W5�Ret�Nh�u�o��ʓ�V���s�������D�ůr�
�2��gVt���9���|��9Xh<n>����*bU�RP�S�q��!�[�D��C����U(���U÷����Ͻ�ELv��z���{��p`����MMt�׬��Z�qj_8к��AX�N���C�A�f+�
b�}�J�n�^�)�SdGގ�����5x�����nf^�F?��i��\R���6���_��ӊȸh���+��·�_���x�A�H&�hV����n�(�/l�ud�)ſ?�� Ȣc��Sj��j��zzz�[����uLѼ��]��)���nd�k<S�ۓ�߻7�3�&���
�VmX6>�-�J�Y��C��ׯξ��M	�����w������zG�Z͋hv~�Pggp���
�{����)*m�9�πp>��� ���Ѿ�׹������K�%�p92���on�L���D�K}�C*����ecÇa.a���ޙ�F���.?�Y\�Y����ĝ����UR�zʗ��d��>8��׻�g�R�-ΒX��l��OW� x몝�U�v~F'a���(p5�*tl�d�x����y��+�ߨ��N"��M��֠���FJd�d�>cv6�VUdnKZ�q�{�X	�LѽB����'�:�����Գ�����S���m,9���C ��f 8�7��0�o�\>���-������ǌ�\�B���a�{%a�۾�a��Թ� �4ek�V]D*�7?LLN>O�^$��s���=�i�u��sJ�����ۖ�7f�J��{�Q��(0�-��n<2��i(eyJ�|q#��.�xy:�Uf����$;�y���O�����m��s�.Ð��y��>���JVcz�3b'����>+fudz8��xD�<:�?��D�@���F�b�����:��s��ݰ�A�+\�f4r�D����������s��%8���s��-Yn>�]��L��E�{�yL�2��GbM����瑃��h�G�~GI�?�  \�ݐM��eVN�

|�0��z@AA����g�(�DQ���9������cc�F�Z�Ω�)NK�)�E@E/ha�
��k��#��?�D_B.g�O��Ij��WwOJ��@�|7d��S���}U���Q7tt�����C��T�A�*�ۋ��}a��:�2	�i4�v+��Տx�V�T�3�#e�	�εi�����q�ړ���z�����\��nS`�v�㠤�D�������Ų�-x�w��N�lA�������|K�������<��;����W5���`��}�������s�qf2eeecGGҴ�4a�B`�o<X	 9�(<�����X�un��l�e�gs��wu��>��J5�����\%��w�J����`���T�MhM������w�gff���ni�MOw��N���rȃ�������]�n�U �K4��<HT�=��#���(����ebb���:_�G!#��n���X�)=#cg�4M�$�?��w��ڄ�����x�ܷ���	��cvV7.��G��K��F��r��-,����]�XYY���RV���tc��0�K{u��������-B�A�ju���x�3쩲���GY�����d�]��:|���sWCv��S�TѮ�+ dzzyc�&x٣�7�*��YӺW�I���h\t�&%� R~�}6���B/c�}� `�����4���?E�54zc�r^�����j����l�:D��S�� �pg�m�Ǐc�=:���y���O%�NT��SS��X�ˁ�RRQ�j�m�}��|�3����Zٛ��Hy������"|4F� 5I��֦-�Ť�6M�6p����>��6� �B<Bm�b	��k�U������P�x(���L\\(���n��2�+a�F���
�mi�۳��]J	7����as����Jh�5UyPhZޘV�?�= @8�G��3�yJ����ذYD~�:����>��2�|�V����5�;~m��z=z�jQ�܋��6_�!d��~�c�:::�؞����y���\;�ֆ�UfM.m�p2��T�I�����w���&������3����b�ى�����R��y��v8�>^�+��۶$bG8-�w&(���2���:��;� Z|�>}��'��pp��
`�%--و�E�'%QS>~����&���M���! ߳~+,<�2�+�K��4��@VR�h�s���_���'b��|� ��Ϡ`�����|�z���hd*)�����aC� ���mJDӊ�===+�g���[&.��OU%ߎs{d�)�}���-������8�����?lz�%��D�A�`��`�XT���O���{�BAQQ�L��j������mfFۤ��3�p����w��B��fL�|�9���
?���K$h�H���x�eT�b�� F�FEE�B���<e`�sw�`H�8/�a�z���m���5|�ry�JLKϰ��nq�\�o�a�+�4�7sqvj�����w����FB@ �?1��!6NG��C@W����+�|�����N��"��e�A�������=F*c]�o]sZ�4���-b�1��4��,@Yz�v+��׌�����ү	~��L7�x-F���2�䦨� ����� Vf��t8_��Y88p�����1�t�8���"Ъ�m�em`��ڹ�x������Ռu9h�UCم/ꍘ��Ϊ[h���V���3��mYs ����t�Q[�����N	��H!Y�wM���U�+͚ &`��3�^ž5�y�!�!��lC��Y��בm���V+C%)��*��ͩ��������l��n< �^	Y	���~�|d�^_�VYE��.��R��\�B��B�Þ���?�l�<�Zn��\�E�@Zt?��6��
{��~��to,7NM�~
ȳj (�x�0OOO�"{o[A������H�M��
���m׭������W~�[]3�<q^���ZDD�h�;�/�F)v>�.����h��"�SB��@�@�$i�\�u����qg��k>>rX�ĺSVa!����r5�]�=Nv������s���\��R��%E���� �D֖ȫwrD�e��J���nB����E�TN�w���5��Q?�|���z�/��������P*�7BF,�A�u�,��wS�o�_@�t���E ZZ_Omy?������4p�zUx����fǆ�m��%#���6f>9�B2=|X�Y�MKn\ ����P�����Ƽ�==r�FT���~�*l�l������`h/�/_�6~�w5σgي���WM$���.}����H�b}����mR����m�,��E��f�6X���|��[��k�	W370=����(���`�tX���3@Հ~=�NII�0��� ʤ��ɝ���v���R���}�=a5�$O[�NՖ4�����؛�+l&_�j�:5!O���OGgf����B��Ê�lj'g�/�%�/ĪG��� �D�:�(�U h�dǌ�)�ix��{��C��ͩ`'�p8l�
2�"��BK �T(�|����*3{b���"3���?ggg�|�I}����䫊����u�4#�)�/~"3�48b@��.�NJ�7f8�k���ܶ�
#昱�b��u�h4�r�^^��I?�gSӎX��=uu���tm��i��/v�Ps_NU��o�Ke��S�|�6�4&˄&nmoWl��,��=���kB��8c��1���6�6�y��2��~�_��̏	��x�+*j��\�L���¢'�B���-��w7���8��v���
w#<�
YNЄ.3��f\�K]	P<�7���ϑ⁴u��4�5��^of�,29�=���T�}55_R�=��av �F� D�w�����8кh��`����؉��5�eX)��ͬ0v(;��#�����c�C��-��{�xR
�H���k(|Fnjc�w��;������Ņۼۮ�ʛdmtMKIn\�(���;��6�)l��Z��L[��zl�x����� 1:v_ |�]3-hY��){Dw�Sϸ�<�큚���t��M���lKE������5Y�+��v�uTb��I.^���0�_��bWztjҀq���N,Ֆ�PFmڂ��֡� ��3`26���k���R��?�Jn&==x����L��b����.�ݲ^#ԤAA�VG��N��\
�+itcc��\m?�&66�+����������N�b~ʕ>�j�L��@Vs�
�S��WDTT�ɡ�Vw�2�}!�6��T$n��b9��?�7{ ɀ�}?Q�
�$�*������LE �����?���G]���$�'�yҖ���WQS#k9M;l�w{T�#��ˋFZZ:�����P�$��C]�Q:��
�`yy|����(#����s�s��}�(�/���0(���LF�Ջ���b�h�+.�eok�]\�]}��c�DF��Ur����L����"�����+.&$��z��H<�Pa�}G��gb"�b�%�f��#2�=�"�d|�3��aκ��U�:|Ř�j�h"�c���Ғ���'ZH���y�˅���+4��X�z�_=�X:v�:���׿|�O�q����&�����F�A_�PR.a�&j�(��A����.?��&���[;�-�ڹ/�*B��:� ����%�.���EX,�l����]惏xƘW����s/1��Qŭ��� �G�sE��m�BZ���>xD�ś� u6������|������.\���s�l�9/���T�����c�o=~hʂ�yj���V��U�jݪ���d@�4˛�t�y��qqqaMmĠo�"��Е�g為�vfCg�}��=0A�1CF0Թ�٨�=��E�C77��Y�2�p9.����ُ::OA��^���a�z�R�(�B������s�Z<�\\�?l��'�}���}P�ψ��;��ի�%�m�Q���b�������+m<h��h04v�5qW"�Mt3#d��k�����VQ���C�C���p��r!���!O3��p���0]�v^�q���ݳJ��`�ط	�r��^��6.�����.�}tw�4�Y��}��̆7�?�5ޥ���!�aC�mhH��df��φ{���{׹�#�����ռ��-~�L�I�_��B�l��R�]�����t�@� }~�Uv�� )a����oM�j�P���s.�����^@�b�f^�I��͞�{��T�ik�i��`�؅cC#*0���KUӛ��Z�hVԮ���������b��7x�݃AZ{8��uˁ��C .����y���ye�烒�O���f�wx���r;>#�G2p(ej�\__'�%i;Tu���{�������(*���*�-������"�Y�H�������� ;bs����6\�W{�0��L�Os���b%�'f5�}��gu�����Lll�p;/��L������_�z��	U�j��֟�hˤBY��v���zVr��%�}n|8��Ҩ�>H�L�g����n�X���+��)_��S~�����߂���!6�^�q�+�Plz1T�	���
��Y~��H�QSS�cj���\���#��� ?�-|_��{&6��`Á<��"�뛺M�<���b�)͋�u�����\~�N�f:���a�임��Ą)9�?�nt?��D�˨�	jJ�6Ͽ�RH\\�rK$�=!v�n0YS�{�0�Jj�O�"&���0�~���ӯ�l�CL)[a�g�����,�p5�ә��^^��E� ����Ιæ$�@=c묘'�4ika����T�o�̌������[#@�]5�s��$�!�=M���fV����T���Q�ئ�W�ܹ���狰eض�H�-��w^)��D6ꇈΗq?	���ee1-o(yz��^BIb����#�_�2��T:��Ԫ;��K��zɕ�;uxH�'��:rNUij�����"�e\���wf�Ó���y��k<8�ɬ������p�!_��St;n��UG�����Ӈ���A,&)q�Ra��b�l�2�!�Y�#`��/��⾸�r�'��3�x�r�����H��)- īE��ؙ��<����LO�ۡ�2KJ��s���0ޟ�>^��B�1/�$p]��A1��n��M�(~lHu���?z�s���p9�eJ�3�t�`��n<� Q$访$�m~
`���)))�W{?珇D�����}/�W����|C�C.����VYY٫K	��� bz���~J9[Q���R�GmMMǶKO$��\K#6�y��W���+����Ҩ�>���ڔR��S����wUz��=PK�D`ve%9 ,�3�%��R���tL}����;�sp�spp@����V�>��M�G�����UY�` ۨih�f���JCC��١KV�J��f����@��5,~i\sJ��i����O�Wq��/�P"9`��pq�������� �+�W�-_;;�o#�g<���/g�4Tç�_�
�*��;."^�J�߱�����AZ2�=����WoOK�1K�k�/���o[��>�g�ڟ��ي}g>]��}��$��ud�>^��ު��p�M?*;��Y�|�軐���<�� �1F��B�џ�ѳ�²����r���G� ]��*HM]x5KM�h�ZM��mᥲ


Ⱥ�
2�ī�F��ws>"	�ˤ��h�ܣ!�}���V2'rwE�����]w��vyJw�.�k���I%�Ǒ,�aB�!�
�?彼�,d�2�~@�]��1�;d.�gO`��D�I��ĕ�4�L�,9՗>���9����\�N�&��h=�<> ��\����ޗ*4��MB����>Ϥ��XZzfa�m��C>V��+uM��!&��������
�����y��A�o�~������A,@r���KJJ���t9�2+�tbƒ\����%�pq'�"��^1�~PUe!_.�Xq]8�� ��� �>5e�;U���Y����̈́�TҌ;8��!؁s�G"jٳ�`,���"�'#"��B4��;n����Q!��{}d�7�_3�;a��&��3+�����ʈS{N�hϒu���d������H4�:;�<�3�g�ѯ�Sn9>t�,r�Ӌ�}!V}l~���x[ś�w�,�!KWǫR�VUZ1Q��ײ�`C�����?H��*�;
xF.�P��[R��Հ��fMKKc�E$�iሄ�5m�ޙMDD�F���� 
 u|d\BBNe%�����N����m�i��;��]ۈ��g ��[V6|&��]	����$�>,W@���z �-�M���Hi����o�2�Ű*dloo���$�}�����Ҍ�4=��E�҇,�m�}�@�w���s4��_	Y��&ؓ��:|�g#���M����}#�u*1�rP3�t#�n{}$KZ
BsQ��������$��u�ܤ�r�O�oA�go�R�ckZ�8�ଚ Pd��&ओ�����rm�k	qت[���;V�q���u�����7ge��-q�6������'bo�K�}6��1�ED���^�Ukv\O_?�r�
b��C�O&�
�S�W�dC3�(�{{yMצs��y�0 ��-4����(g��E�D�*&6-1���d����H<�67 pfm�W�._��d?��h2�=1#m0]İ)��֦�tu�[:���� 7mr�w�9��﬈�����怆�).��OL|���y�j�|��?6b�.	�-s'�-Y<<��	�մ_�Ud^��mE����i�#�RWg1���y��l_�حlh?��F�$'cϊl�FC�Q��]�b���Ғ�L�(l2bW�&�Q���=lb�X�_��`o7&-*J���rPnٯ��s}R�hr{�'i�SUs�[5M�|����(��.��6kg��;P�gd^�`�Qat��c�H�Vxr����(��N�r�����)��3��-V����
;T)�{#追bf������n9�!+�jZ�\�B�y;���22A��'�{�|�*��������6QTr"��]H=@���(0�����6U3n����?ޗ#߁Iw4��V �#�P� ����O}y�ԍs
��w덄4�ձ�[�'���DJ��i*~}��{a�b�z��T�jq�0k����ݡ�QI�{��V���kf���R?���M�%���1�xx*�Qg?߂������܍��~hb��� �5R�c˪��VF*��|��#��Nf�@|FFFy��"]��~�({��sz]��>��?دbٟ{�<��"6���')�P����K�����EE$AQp��P�x�����\�d�&��v�!��g�m_=A��F/]�7�����W#e~�9�ҽ�����[�J1A[z�� �������T���f���I�ܗ��j��k�Z$`!K����]
7q�ۜ�?��Ԥ7��_Eyߠ�ߍ�/4��	i�4��"Nym��u��W�d7����$7��m�l@�B��~��?Q��ؼ�g�վ�e�V�׷o�"]�܆BJ�ǰ�W����4<���'��o	o����q#�8���55��������fϻ'���j@MSn|R���K�[���&��hh��f�f���զ���4��LՊh_
.����w?o�9�w �#�j��&�Sx�1�BKw;������f:�w2�=mi�Z�޷���q��B_uG�I�T���=� �Ζ�������Ξ��``���l�-ED-Q�~�%;H����
aJ��4d�	Rp��^,�un#e0�Ve�E��z�A�x�q�z**��߿����a߾�p�r`o�n~�U��<?�7�[,(x��_���Zq����F�I��Or?+t~�����u�|l��'��O#�F9~'kg��C,�ꋼ<��0��_/�g��T���rmE�]qKGdI}/E�ϧ���H��G������Pm�kk�"�����kO�ߔ��
c�`0�
ȟ"�0�ͨ�961���hV_}.�$������^�c����C,��� 2����[������5�M���6�%��%N��$%q%��$��� �qܛ~�%h�$��iq�TVV��Ɉp�$�����Jr%C[�*���Ύ����oe��{�ju#s�s�bSs��.�c��A�B�e��~��.�UCSs�l{<�l��:ӚR��X�ԩ� ��H�k^��c"�����[^��7�N��+=0�OÓ�I�f;qkn`�K_��,+���u��󊉅mo[�b�j �����f� ��B��N�}���� ��q�kc�bbcc3[Z�o����30sS����
��)��K��U��g�c~兓9��o25\:��������tp�2����**)��?~M�-q�9�b�:��5�hat��
�P����9�SSe<=��m-�?��)>��Ȉ���e�t����ذ�c�{��>;�g����.ѯQ�E����yZ�f��]g�
B|��9H��L��o�π�&C����bb��߃��������6�R6r>77Ǥ0s�F�&\J�R���$6���Z����\)���d�aC��ӑ�P҇(���7s����T
0!��4%s'`5<�~����/��/�v)�3/�����=?�ۛ�Q��dm�74�`���㹎_C�J�h_�WW\�������wdj�EAv7��!}Q{�����'Y�{Z�����{��_��JN^>�8=���:�8���/��vIdp`l�$>�!^z�ط���D�6��Lo��3?�@���������ׁ�����X�K'dI���!z@��vAF]w�#abk�\u'K	����^vkMX6{>Lȕ�x2;c�	F�Qō\��]�f4�*S���cjz��b��kɖ�C������ϼ�o����� 
 -1c����B�0� �yW;��wJIp�@@^��J&!3Ǟ�0{��������]}ơ���64���kD^�^/���d�fߟ�-T��x����Kw�1=�'b:�;��弼�i�.�>�l�/K+�����-md�2����ڱ��M�p�p��^d�!���T�SPP�2EmR�|6�,�p˳��Z��������d�E;�k�u��1b�!v{�ʷsJ2. �VvώR����V�>��5$�4��e�FY�׍o*�� ..0��>yw�f�dr6�DZH�DҬl ���re�7�*^�W�P��᱆Z6�� %�J��-� $���;�K���:�����������iy�\�V������{]����-$�֋U%�b�aU�q�B��UU�A$��]2T223Xg���8Zr8BhڮfI���HQAO�s�8�YS�^P���<��Ԑ��=���6´T>�X��w ��Yϭ|��:E����|��YV��3 � ��5l`O�`�k1�����@��g���h�~M"�� }_%�n<ܸ��C���+p ���+�S�{K%���*4�466V�{�}y�n��\I	��|����Q��(��X��+�����������A��D��n~^�����2��ǀ���O�W������^]��=���2�Hp!~�6Wm�p�I�}�<~���s�S/o�c�	�=��f�KS��Դ.�����%���5&���&�6�hѬY����?�+���#㚝+��qd�n�'��< �#���d�e{M�2/�Kj���ဦ�-�9�q����7���55᪝7�ebuq���{���P�ұ�{rrB[ 4�
���w5;��="���e��ݹ�ɰ�!��e����=7��� ;P��/dk �i[[c�6�Т�.��w�Dtz�A
������C�����)�B�,QNNOV�*k<�t���eQ��DO#���*���;�Z-f%e�i�%������9Q�g�ٞ ��6aߕ���Ybkt?���v�������Rw��>��jQ�%n9Y�{t����7���M�YM����6՞H!��`�^��n�/:�w��J=��kr�K���|�~aj*�(�ۃ�<�EE��*�!l�+]k��Y�Տ����C�K-�vZ���uu�Z�s>�����ۗ���K��lO8-���Մ��jX�4Q��c�hAw�:%�+dV5s��f
D�����F��fΎ=?W��sÍ�T�q����g�z_5ha;��K��>N�p+"xǄs�b�Ҿ[� #]Yxӭqtt�	(T����jj�ep��Y��JNiM�NoWm�6��n�i��XY���봭{=��8�w��s-D�O7����I�"x����^4�VM]��L`����R�444�o�R�; I��+;}S�JN�P��	��?���.(,�<�.x�'�S���N�A�0�S�+��T���A�`6�m奻��o��pՁ��&���ٿ�q<�7�O(�)���.Ѫ��JQ��B����S]�mlLC[�A��3$��(�6�Mx���ӛ�����O��A}��y��ރ��wP�,[ܯOb��j���h�E\6���Rp٦ �n�=��=_��6�tv柝�S32�x�F咊sV��S;u�.!�5��S* �A��v������Qԕ��mq�K���6y(�df��Top��-U���UI[�3�u�9jaaa�vv�����rÐ���\\��������CdI��N�7��k��on��3���;³�����7���]|C�����2��P�,U����_�����:���͵h�֖��G\� �ֻ��i�EEX9��3������TT�䮬���w𝔹++I��_dd�, ��Ȅ]��t�@�>b}��iVE���Ń�Σk�c����۷���W@�X98`�e�C�c��gH��P�����j�l��ν���'E�loo���'��D�J^^��_�2��TYii<=}���y;�+�B4�Wi7�k���@0U��b�Ҡ�ᯝ�g�������S�6N0�J��o �r�TE�m���=��殑�e���zݏ�wS�Pk�G�n)����D�a�����-��꾷a��A�E��SB�FR⡻;�K@@:�S�FZ��C��w���oƑqn<�9k�uŎu*�.��+�����I]�YXX���7�s���qt����$������E'd�ۯ6'�+d����u���E���?s3|�Nslg�Ư���,o����{dWk��k�Lu���7��555�Y��Q��(�P�xtB�Ռ�9�������
�(�S�{X��>O���?��(���86<�]��*`9���G��Y���1(�}k���=�;�ׯwo���`@��g��������QW1������ug?C	q��*A*�����Z�ۻ�mfo_���̀�R9�,���Zvi�W��H��;���zr�P����CG E��=����Ǫ���qlt�
%u��V���ޣ��̋X#vK�\e�s��Ж�fT�%����T!�m���\<��N^�;���0ҭS�R4����,,-��U�m�ڟ���ř�e�̷������属-��PR���c>]Y]��6T�lVM*����՜s�ʊP3�Hg (����8�b�ҥt��%u7,D�V{%#����sk���jP��ݫ�Z���ߜt%k�Y>ZukIqu�S�-.EiY��d333��<1�mlk#��V��P�s�PqFD4����`�A��t��9=`�^��SV�Z]m���d|������@�!���ڛ3�ۧ��؍�[[Tbbb��@��~A����3d���-6�[?N���gpX��L���MK#6��+�.���ɉ�9�+J��ۛC?8�_-�\�޴�%)-�S�����cc������j�m�,Z���C��`�7��Lv(.x��FpQ4L�(�n'gg��{���r���8
�`*>>�9C��/gj�:|fQQQ�7{3e���g#i8�e��|�����U�p��]�X��~A�Ni�a�%��#l����f��;>6�ɡG��7\�ʾ��p�8Tc�j����ݨ�����O|&��.:U�}��Hu���ܷ��lnY��Q3i��ɠ���!Q���Ekǐ�z�ذ`
K�W*�j׍}7�B�����{�/��r�`�W�3����,?yN��8^����'�]����=��ֆ֫�R�֮}V�""�>�������Ņy��lᒽ��k�/X@2Ì�Oh�MT�8Y��Ʊ`&��0��]���v�S�D�J7*ӿUZ�U������"k�Xސ�lSE��ܪ�/��R�y���RSX<n��05?k`��v�r�P_��F*�D^**,Ċ�J�Ɯ;��{�5����W�;��_#|+߁�K�~��l����+0&EMO�s	��U~�ӑ�g��T[��eϬ˗�^y{��^�k���S��n�@RM��UP��-3@��:�L�z���rtu�A�R$j�- &	�s*���Ɋ��&п��88@nǩ���8n���}B�n�9�?//�ܕ���h�����o��ϡ��!3��Î�]���艌�oܑbA���c����"�Z8
��+)aRŇ飯�>�q���o�C����k9�I/&m�/-��o��'���~m^�;��}󗂔�)�#S� g�+
�ȵ�="�*RzA���^����JF�i0�B�m�C���������8ϖ%Bs�dQ��ؔ��(u�|Iy��OO�,�s���|���E2$]]��ي�V� ���姞+!��r�ͽ��7J�'/�;`+�����2�EMH�uU+��o��T��<B��m:R-������*.���K>־4Q������N���	II�@vT-��Ny�#�m��O�g��558	�Y(�8��3権�8��u �ѧ�:�#]��v��AGgy�Y�500@������А<�A���i�̸�aǷ��9�U�CujYhU�sn��C-r}��תj �BBB���x�!`���B1|֌�W�_�ް�M���z�Z�f�&�z"��k�矼UU��!��`p72�w1e��+E<�j��# ��Ny�B���+�Y�Q�]~@�������� L	���y��2�;Ǧ�CD��g#��ӨV.�L ��*%5�C{Z1��CUE���� )���V�߆5gD��tTF�RMaiupO��L�8�*�Ə�(�Bݴ,Q&���(ny�1|ձ\N����.��Y��A),=-�z-�Į�E�pPl,���jY[[<}���¼ee#���
\�_�z���\:P���`
��r}jVV�J���{ը�]=��CA�I��M��ll���?��	�@�P[]����16~~شM�#I��А:��o��,)44�r�KWp��痵}� ���w>@w�U��d��_�}rr2J����;?�V�KQ�7�����h��kRz�	y�IҔ�)����0:rK�>�O��:�UQ�>pkɉ�]?^�%���%r�\ԋW�9���Z�w�0����*�@������8u��c"���H-�c�����I�)��bb����xl���\G�B�e��v:+�2�!B�''X(�Up_�nf���R|+��QP@��4������� ��vɼc��rkq�;��b}�b���?�~�{�Ԅ���R�!%I_3w����o�%ɶ��/45G�,�c�M��D&�,:&�s�읩)<P�&&&�h�/A����i8����g���������VH ��k��B:�1 �����������IN��k�E5���c�H��q۷����4�V��VU���ч�����q@H���T��y�������q�5��-��cN/`w�=��7!t�|s�4����=�L��t�o�����%{,����n����\`>@w9f:\Tȅ®��<�|>����O�rJ/��Wk�j�������s�7�JJJ_�^������yK���	�[�����w7$��1,-Բ]��j�ͤ�����rZZHD��\,-���:�����deb��\�?Ivh��� ʄ��hH�36��S]��$�e?ػ�i��|��7yY�Ka����t���;Z3�k�q݂��k���Ύ��WH@;^�1�{~�4��"�Y���Y.��@Bf��[��������O��� �F}:�F��W���$1��W/nօf��	a�L���8�,_�����Z��~]����Ibh�^��}q5�S�P|�{_�K����ll}d�K�P�~�[�XR� �"�T�)�#���IZ_�G��a))a�]��Z?JY�s�/1��S�D�����#���T /(��ZgY;�Z �w+����K���u[��_׼�5�ꩬ��tx�������o�l�/Wƿ%��Uʓ�Sh�
��OJJʓ���4��O:��0 ����	�GN� �EPl�ywV�ɳ$�u��k��M?r��Dd�+�����se�fQ�~��:#�[��M~<h���I���>����R5��~|a!����i�q��Kc�&Q ��#*\��:�(s�^��M�E�������}\�f�š��DR � -"��r��ޙ��6�9�'�Z���!��r��ɠJ�uޏ#�!n^޼ϟ��]���D!.E�����P���;���A���i�R�B[\Y�&+$lx��n�tS:���g��i39��V�;�����+X��۷���l��򟪻}�Ԥ��^S)}���6K��s%gZ"��\���� �ﴁ<�%�*�"�"E$��~e<��x&�o�����N`�CXj�߰��;>A�+�ҵ���+k�ɜ�>)���6�t�9Kf��Z���9vh�tP\ZZ8C����W���ϣ߮^N�ec^mz>�W�ۓ#t{֕w���^^�<<4͵��%�����)�G�=ɀ���g7j��K��Y	�~���չ����J�:�=`j0����a���۸�̈"�L
�3��
Nxx�@��Ij�=O�766�YG���	��(�"`��&|jJ���I�,	��,8DEc��*�23��Q
������p�������~��Z���r坴��:��s��N��KL�F�3m������]!��.���"��'��[%��*t����(.MSm����g�XC&��#�^�	DT��#��v�Cy��@� �n�Iސѯ,5�I�-���� L�KL\1�!���/�� �x��%}A	�	��������M]�|��Jz�,�=��ߵ�-˱����ZZ@���Κ��tQr�Qq�7��fWy%Q�+W�ik%����e���}qس_��0h�z�J)�Y�DcՎk��{���Yf��u���wՄKvV	��'C�DD���0�dGu��޾3����\��{~���o��D�4%��|�(���[��DP�|y���q|�g�UD�b淛�T��|�-	0�7i��9W �_:}:u~���g���Do��Ѽ/_��y"�I��E�(�`�~ m�����TTU����S�Y�\L�	���x�T��4�U�)!��B&�ֱ�WT�Y%A�#L������o�`�^�mf���f�9�y'�o�8�����!��������JEpC?}N����o6(���!����	3��vd��N�O�����EQ��4�[U<К���<4�7$��4Xj����֪��|2=-P�h̙(42��'J��q:;:v8���s��sW���&�ۙ|�!�;�����F�{Y��B\��K��}�'�2��5S�ߵ���&��ЩbyyT�
Pl����jSd�s����@�xq//]q����q��ɨsIձ�R�3�Ur4D�*���&��4�x�!~׽�;���KK������\ �񤢢���.t�r4�W��b�;r�w�CI))���ؠ��t8�+O>��f�T�F������䚫c�j�D���TM�q�A<�Z�w�>r�2NA����|�Q�3P �걆0�T!�`z��о�9`f:idU��9U�Kף�	�q3*|I���I���n�F����xC�/���7Y}C�/�R�j������v�5x6ǲ���s%���Q@<��I�J|Ս��#����'�g >��66�4������7i2O�Zae7.n�Sĵ�SR�[P�yc&Cɽ��[A��PJ%W ߽�0���bM�]C�CP0D$P捂��R�s�P�`ww7!9y�[{4�����g��GҕI�Ʒ}��UUW��Ҽ��A���|�Ǻ~Xh9ݩ�<��;&�	��/��z�/<�56�&��M�5����Z&^ӒٵW�]9���8���:���l"�e��F#�+'0�u$.�j�A��o.0��$>lQf8�����43~��g�� �sѣl�XsflX�챢�8����rl�we��c D{�������j����͗\3�Ӕ�(#����������VS�u*���8S �yq����hQ�r�
 b_��"�����8C�K�%{�J������X�����+nv��*�r"@Ct<\(H�h4�۪�3�f����Q�i>�݈����>��ʳ���逸��Oן�7w(;�?������10jV>�-���[�X"'%}?�R�Bۈ��~��H�/��{���Ó�!B5/"n[[P7���	� )��ޥ����qG��/<:�4ssJ\dx\�֌��ܝ[�ve��?���r+,Q8�O�L~�����-�Sg3礥���?&&�r'ڪH��,P�H_�����.^_Ù���R����Rz[�4������м�a�A�l��<�ܮ��^��ܕ���[��=0@�v$###rl�[�:z�<��%q�e�ܚ�*������QB�UCA��٤_ثl��]]XHk�Ҧ#��Cpv�le\�l�kׅ����䡼������z��OS_����_S�k�&`Thl5����+���m���Dsh�69o㲤�F�ӳN*�k��JCC3��"�Ðe�i�N�w��,�����4h��j�V6iқ����=���P�Y�R^>*o�C�A�+EE�i���]��qJ<12/�5�d^�2��E�/q��qzܗZZ�Bs=��g�r��a�S�%�$t&�dd�WVↇ� h�����2
>,��������k7̴����(~�
jOn˫�m:=�B��swu�H��Iނ�J��Gqd8^~@����,A�����ڍp�=Wx�С_5���	pB�Ȉ4p[���[�s�	���_��\Y����m�������(�v� &�[tKN�=���]C��U	r�UKl���o)�8z��������B4�eЩ��6��F3T����	 �n�~wN#�%w��}��g=W9���s)8C-�sM��t��n =L'��[`Ʊ�i�"�#onn6��&��G*�!~:�]`<99���]�m��}\4ĉ�Ũ�[��mEs��\Cdz-n�A���4
�DcNH�f̣;%��P�lT��c1����5��D�z�;��i��~�[�&222����ɾT��AcMAժԓpt<�ӊܞOM�1W�l'i3P�5�8�8
HZ6�¸��}+�FI�h��&J<N'�(|��u9F(��S";�r��!o8e*l���BzҪ������x�Z&�f'���2�-l�zk��+��25�t>��Szzz�����@�����Sd�����ܓ���I�����W�@��n˝
%Xl�.}�"s���p��'���e�����,�C����H*N.��Ag4|-: w"�Q̰��#�R �4�47�|Y
����E+3�����BЬ�637׽~L�۾`c��Q�Y��H4t���Bĺ�:B
�㤈��2��=��Xw��SSp��3�Ҷ�g�E5}�k�&:�����e%%�?[��t'Ё��nVۯ�^��.lHc��T13vrv~Vj���.p�&th3�aԱ��$�Edu"b������ޝ$	\�n_l4���V���v�z�|�8�X��=�4b�N��ZN�� �@=�P�콅���U ���krss��cqo66L������N��8MmiV���g+d��F>Գ��w����eJ]ޛ);����ck�|�f��������ff�C~��t��m�d��Z�^RES,M�}�GGq��N����/Q�?��x���*��Y1Ǩ|����b��Bn�fC}���X\�n����f����46�Bz���u���5��u�U������5�^k�� ��D�kvi��X����>#�\�x�T��a��IS�~D�V+�W����闢�"y����tt��;DT�x�ޞ7%��X9�+e[��%<�M<-ԏ����`FqY�߯��a+++܊u���їz�ys�/b4���T޾��"`c�e}�uǧV6S�'1.$i浴�T�:"��G���� ˁo��f��F���Z��F��>�&���E�n !�� $�p��p�5��*����7���s9R2��֗BP �ց!��a���j��YLi^/�.c�:>J�.Hل����W~~����	1�
�=I6�q�;|�+��ᯜ�c��>�>�{�RR�Q�gM�ީQ!�C���gTe%�������֎3�e���  u�]�0��얊�o^~�x���_�T�5�+�g
¾M�_�~��q��Od��UhF�Y��	�˔m�fJBI��}�ۈ��� XZar@�8�E�xR�SW���=����u&����ju�ww�rJ�N-D�[L�CJJطo�)y��#� ;^��W� eSM�oo?�V 9���,U�@@�N��-��^��g%I�?p{�� "���?�%7�-��6�b@�5 ��A �.sa��8Զ*�Ȅ������5�E����<�$|�x�P#]5b�����jM�/T8~�����9���}xx(C�+����)��6���XyE�ZadA	[9�e�'�7s�Ʉ�R�I_,�Cʇ��2jj�y�J3�}Ts'�,-w���4$�R����	�d�ۗ�W�����`?0�.X����J�{(��W�GZTdd���	�씐�R�'�A�r���{~.Ãega :G�����[EQf�V�|=���P���6��Bf||�����MSI�����e/_�������&m�di����7.��n��TԚ\D��i$@�D<2i����h,9r�"�ꦖ��t!��x�#��s33 Uh�`rj���T�i��}���Ԓ5.��6o�����H:�R���@�?�G>H�W��}q�|��w��w���t���y���|xV���9�I��,- �*'���ݎ',W*�?O� .�Di������@Mv9����7�%����laa�EA,UAZ���Hc�9"F#<8(��d�	mل�㻵pǈ�������T��Nm�����@$��j$@��!��>b����55�[%����Xq�bk)�Э�gԸ�#N�s��,���f$ԒS3Ԟ.}�7��k>__N$����U�貁�.�ׅ�b�Ap��.g�B�|w勋�?��ϾD
��HWz1��,�{vh(�l��ۦ\Y0f��ݐJe[�������� ����/!�V�Rg&������I� l��ի�߀�	�8a"�p�iJQ�3���&�f}�9V�)+G}!�����#����������:ؑ϶P�Qۍ)�F=H<iy���(�mF Dm�/�Ό��`
9wLf�+��c����Tjp�};��e�-P.-��[���)�r��T�͝�}�����I�j�-��u���k�����K���D����{�eUU�:���%@s�=[qH�����k�}}�T�m��iQWS�� =O����o55��E /���7uhR�
��� �,g�8����8�_������,�k	m2Ҵ�KY�Z8��	�2"��'�%fw�)x����_��V����W����^it\"�+���zB���������п���0r���J��C�*�Ғ�@3IQJ����@פ�_���O�j��b&D�)� �y�"�qŃ�jRb�י����RFBy�܄⃨b5I�p��������104�C�����������C��i�hUG����qP�5�"iq?
1o)��N�$�,�����ll��%�hfq��Ue �Cf��pFӒ#<<|�q�Ă<�����$Y�=�<-&�����5�Q������\�}O��e�7`n���#t�XR&#���T��Á���J�����C�ex5�����ZZd%�-��gZ�!'''4��#������95{�lN�9�a��٭f'�/L�-7~��[������FHV��|�������f2�܅m"�d�&=�MSV���`\����͗u%h��^q\�����دξ�װ�(y���[_�9����{��1�I���`�a;;�McsK''l��W�kX7 `�r�V➞>WA��)�If<��>�iii����2�4U�e��H��1��-צ��Wu^^�<�1<���1�	b��۬O��6�l�}�>OX��X�x���/�^>��<#�E����^�����꽻��{_�3�H^�Yn ,�6~�g^����sU)>�%�J

�3�GGG}3eZ*����`���(�o�U���������Ē{q���<���j�f��F�M����i�Ҳ2�eU����]\$S#�6�/�L�||HA�V�d�C�K��i�q��m�Ad��^ѹf�tEIsy��4I��	Í����+�_QCt�I�>:��!ꫛ�7�rs㵖��(3�sku�z�[ww�%;�7�� �O|_��9�թ8�×�����a�d�-ll�]Ї*2�U��>��HS��%I�UF.R����w�4u!.���!�?J�-~�C'��K�gaa�O�����߿���T@*ּ����0k����rRt8!�\v�x�3��<�_�]�@~��V_MMM�(+�����|���t65�.{��-#cԤ��ν+��(��|:�j3_+���@8$܊x��)n�:ʦ���2 ��233�}}}�e#׷�ԧO~���R3윔��#Fy�4�GU04`��NMo�� ��;��'�i6�|d:�����r���$�_X�A�)�4*��8Runl�܆e�����*&G鋣����C����0�S�ʪ�U�	�9���K����r��O}^M�j�U
*�RÍO[q�/H6��
]�
*e���iR�k���r+�:p�tL�j����}iI�gˠ�̬V��W+u2����f�m��{k��X<(ka�-&����-'V�������puU�J++5]�y�04�n�V9Z[3��n�$�=	F�B��z��S}�	�~2u����W7�h�H`�e: %ۯ�����3!�Q"��P��F�NS兾�,0~��=ɇ^��}�4�i����kt����`�*�� �B3m+��KAA!~1P&�"�v�Q�Eߧ��7��ܿX	*�E���F��|=a�gF�ګk��}K�Q���ԇX���y�+gzܮ\�0��6�<�f"�eV��m>�O�{�MN`��,�
rs%&p�i����#��A��������XD2����Tk4�gX�b�~LI*�e���5[�� �qu�G^Mu�50q^8Yg0"��5�[��
�����-<��v�Y'�:�����0O[k,�6��j�Nu)*�'���N*ޞ����8WUֽn�/�����(�r��mͼ��sh��i�4<�g�`�h�{r�?��Tز���؛�U�oUT�L�6��Ĉ3ss��E�U����������o�tX�q��n/{�����9j������
\$���S����/����9�}7��K��96vi�3��v���/�Lԇp{,[ˈ�ƌ#�á��h�ρ�˲��� MԭQ��(�V[QƮ��&߶?������A3Q�'^�+����1���7'��1N�o��ճ�+��2����4Y�AV0��m;� O[����SJL_�u�32HA���L�?�o=���D�^�&�F�Yo�����d�IYWO���/ ��y�󍎟�N��;a2�kX�� ϶t��������Z��x��X%4�7_s���%]c��/0]m#�kL1�%)^�����gez��b!&gH��nCK���!�ԏ��je��
#z 5���#G�&,� �׳��G/��/|y�Tp��n��k��s$#6���$���<�.�bl���,����k6M�S�/��-����^���eƜ�o���	�^�WI�w=1)q�a��XݕG��qS;ϕ\���Qebd��m]�aƗM� �-�iw��������<�B�@�S�P�-?;����T��U\^i�\�̸�G��++��+U�K����h�iL�r���p�-Z[[�;f�-���"�wL����(ur�4�Z?^�Y8�Z`�N�3�O�}�LϽZh��_���<.�M��Z�Q����D��ܭ"�)�z��(���t�3�+�XZZ&$'�V�֑-�|�;y�O|y�������U/`l[�Ưe9���%��c�܉*'� ����G�Q��t���XD�:�I���o�����v��R*���ؗ�X�i��%vvV]�z��R�s���U$��������i��-��W�����h�@� =���k�V#���
 j�┅RSeUm(����韈�tOA���������T��U�Dk����WRΪ�G��*6v�����lT� ɳ���y����M�e�D(��*T�hd���Ţ~/Y{���t�<zh/�H�`~�21	ɚSU�'��)�JP@(����3%JJI�s?�19*_ι�T�n/i��2�%Sނ63�@��(M�����S���3�tM[k�Y��D����q8A����I��P[`�`��H���XY5ˉ\���؁���)� ~���n���2Jt�˲���S�{�Ղ��D��b�|9�5�o�oZ8�p�����d��o`��ؑ��W���G��� ӗe4��Z�F�9X	ӈh)�ˑ��FB���лIQ*^{Bc�P�4��s?m��i��k4S�@����Z��T���b�:�.f�m�g�Oګ��]F����y���Kp3����P�|b�!BCP2��X���g+
~�ω��>5o&=���Y��I�+��zC[������p��O���oX������]PP�E>>9�zF���t����~��Z\>��5��cm��ZUH���?�4\&������v:*�Rn����k�Q���w΄�)���,�F���𐽚<b
���l���Q#�đ��U�ԃ��Ы���]Ϳ�7��ybU�|q���7��p*����e7����J��dx��D�4��חvA N����ݥ?��o�����e�K��w���t��pQyP
�璘7�	�,�R;�,���d(NZ���"О}�/T�P�?�3H���f�u9]9��X�Ntrv68��7k�X�m#�lY!\��\-#�F��O�J�W�U��=��v�A�B�;s�.̀�7ͩ��ޞ���t��<f3���z|�8:���B�����x� �_S2%F����Y/��r�C�����P�_��뫜5l&ggǕ�3��1�����obbbaa�t~s�qشmD?Ԥ�c�"
Wm�2p��L�^�×�l���7���*M^��(��s�-F	,��E3����g�V�NN8lm�T-���w��(�ӻ���/[(���)D�1�����T�1߭��D�f���yC���
܇`��d�Q[��5?~1���"ֹA�jm���T�YYB�-�l�/��-{m]�'�}�VV(����í�k�~�12'M�A��0
�h��Bk�}���~~8N�Z����⇋3[���X�n{�����b)C�K�1���j6��yS�Fu�4l30���*$<�f<n~7�_�#L��;u@���H�9��*�~:��Ň�����%b�������f�5,�5-OO�F�Hy���>�x�'��u�q��P�߉�MA5������H5���r��_�cޙ5�F 
1O�t��� ������j;wT!�v[n`{Z{ҵ�,}%%E�ݧO����m~-��۷1�.��w�9t�9��*YNurv�K����jV�k��X��T�U%c��j �p{�z�#ҩ����Ήm�r�)|Rx҃��p{��~���݊��ʒ����ů*��}�N/��׺�N(Ј��HHE����;[����i����Ɗ4Cc1��"�O2r�{䝐邑�F�D}܂ہ���#�,���n��BBn~4x���e��e\]]��=�h7z�����V;5D�4/�<yO�?��:�'��T6� �2�NNn<�W�&5Qu�5��D�Eg2�P�F+gfvV&�f�������x:��
�onf�"(��5&
l���ꖂ�׆���ߪ�)(���Kʩ�w��/���,��݉3�W��CT5W���gy��7�\�>��EFg
8#�eH�f/�L��}�Ŕ�?y�E���f/��ۧ���<锲�o|�ch��L� J�^�2rq��7.6:��OZ��T�������c���ۓ�����On�zƪ8-sG���_Q��x����Y�?c��K@����Ωoh	ѪGƺ$Jq�8�%�z��$��'��WP@GDD�j���u�������]�M?Qg����|�0(6���>��l�� zQ/�~TQ
X�5�~�=�����(�v�5�� Zm�L�In�3#���Ů_����8K�0F��5���Q�䬦7�Sރ��i����oŉ��F<��q�*�:�Ö�vkџ��jm)m2���hT�~����`�o�~��k�fRT���w��^�:�<��C�L�f��!��E�~>4OI�Ɩ⓵��d�x-c2���zrs��w�-���{<�ق���(,d� ׉������x1�o��q�$멈��?d�P�퇆�|~�.v�P�����Y���`~Qۍy���$�zF̈���Ϧ��
l��u*ZZ@��f���N*����a<���(�Z��o������4��,�X��c�����i���Ӧ���z��+Ր�Оw�o ����B�h��H���2}�g��W��4F2W��3<<��R	#����e����v�Ҹ|H#bǿ����&��BGrV*1)��[Q�)����k%��
4D�KQ(F~�b�n���߼W�7���t��?�0b_�	/gYiދ]th�z�L@���e�s�>�Qj�DI�¢p�l�I��CE`������2�T&� �������g������9�0ho+r�u�Y���l��.�ަ�>0�r܏�m��j����M��^2�LI�:��T��U6в1�5U2|0}�v�SA�s���vFT�Q@�ڇ�	`$�C�����'����w�Yf���A�ЪRZlF��J����ᚡx��d�E�Qns��D\�U}�Ѳ�<?[�i���@o^��g	�����8"������)�c��w<8��&��{F2O]_���4�x�G�̉�x��<�n��_C^��X�k��6��*�k���6]�����̞ɚ�u���?�U
+��2Z��L��_:���U�G�|���vr�)2�c�XC��Q���Ι��߳߿����|�K���_k��"K��l}�|����qn�s~$I��{�����Xr��G>�d�%n2���,����4�<|���)����J��c<�ZFn�Z*��p1S����Z��%�1�GtDɥ=x4��(ꠓ���'I�M��Mӭy׼~;M�d���>�_.eL�q�E��|q_��m=����!Kl�D�L_�1:0W#7�A����sz�x�L��������X �+�8�Ͱ��;�#Ńlgk�sw��@L8g:P�aJD����dΣ��*���dC��}��=lg1f	�׆�-��A�	�������b�ʸZ�W��#=i���N��V�g/)/GC@@��Iw��G�8�>� V�>>�w���%�U$V�ݬb���k{V�h2���%�码�y��F;q� ���X�[&b����}�F�}��m�"�T�E�-�'�qq�iԫ������jd%�m2�	+�1�g�@�5�:Hͯq�{�7Q��hh�n�����8e ��~�����"���ԞjvV���
�Pk��F�I 	���vI���9|��y~�!쉓�L��v0���nT��.�mn
Cv��*!"A��ك��Nt�cY"Q��a�ጭ�#�{��^�	1l*���1׳��v��Up��ܡ��]5-{�]4���1.zII��޼Y�-��<����I~'���J<C�p�Jhz�
��`.���ҳ�Vd�ӟZ)&�98kv�q~h�G�N1��157��E�X�K�P�N����N�j#�����#0_�g^4��P#��iqͲ�/�����"mr�01��s%����"`���_��V�Q�m��5G��K������F+ѝ�X���vv2JJ���狳у;j�-�o��[0Up�NG���(s�|���-�C+##�G�����4�������Y�f�`h�&�a�ͤtl������y##<�)�s�l[�#>25�s�ۼ��D2�����
(�#�6���b�՘a�
(*��jgv4d��8����A�q�ܲ���������?.���\e�I�:zVV__ߥ�J��#���\�r� |�H�k,x`k.W�1�x9~,.'f��o�=�?f�Lˇ��w�L6����2^�}������s~|< ���u�g12%��i�X�u�;.��w�J�l!���+U� e�����q�\�h��ŏ[[����>�t��"K��D�_*-eX+s���]�d��ϙ`�3�5�:՛����c�ǘ�����k�q��,�=֡�����!y����%&r��P`Da�'L�L��-�v	�TS������8����|�AB+�*)�lI��w=��'>���@�ro*:��~����)���);�8/��)�n�Z�iK`r8->ԋ`]Y9�:��+���=���r���-���*�ꥼ�ֲ�Ԕ'��sz���8����2"N	�`�n|VV���M��!%�7g*��{�5���� ���9,��R�P��z���7���Y8������> acӈeAǦuc������V�YPص��O��n_L�mBg9�����TW�5f'��,��ᡑ���-�d��������1C�����c��[��rƮZWhƮ�`�蒝����)���D�juT���"�ņ�SdXh�\�%[�vOm�c���d_�-6���,;��h.��H�i��Hۀ�KMM���Sh%6(��̬ӆ��Ɛ�B��"���ݼ�JV���9�>o��C���Zڷ�u\#�+Lӕ��׀-:~���eՄp�ֺ��w����	&HW�G�pc��ũT/*
ʟM6"h���HRE��ʹ"��\���T�����#����\;Dѫ�_�7G)u��P��0�"5n�4�� �`������@o؍�,R�s��u���f1���A�,l�袈W'��]��Y�?b���,��j��)��c��1#��҃�HN.|������oB\�~w��q��ᆮ���$��Ze��=�L�unYD�*���e +��]�O<�e֯�dBj����>}
�y�i�pf�m�۽}������><�\�MdMhQ�z� �@�b�,�(�� �ê�%��s999)��D@;U.��13�lr��jLU���IH�;��>+փ���H$ħU���B�V[S�*�0�Q�^�ĒvڜLF��I�O��X�C��gg�	Ѻv]����d>c3&Ev��K �$|��C+�2p����^�v��?�g�o�L���<)<a��S��x���9llU�I$w5
��Ɍ?��u��Q����*>��J�������Y�8��*d��Ԫ��7ݠ��5��L���
M��6��{-/l��W"@��00�aa&�����貿�N����ϳ�~��&��b�f�����:}/�	Ϊ�7��5IO�I���xrgh�kc�:�=���N�$�/eha�����-�`�!�!�f�kD�0f5��i��J�7y�!%S�[�����J<-�7�_��W��F���)���5�:�.�A����NX|t!C�f��<a��OU��p?m嚯�2I����N$
)�i�&=�����m"�{>��^֕��'�5��#h�nU ��'8�)J{���s5W�ø���c������*z��o�3L�8���_;�����1�0���#��(>��\!0^��*)�V}�z����<��8&����Dl�
�VU!�f�tܸj�r�Q��#}
�`0��joCg�>����?䞜�̙���B�U$p�f�'%'�MT���G1�X��p�9�+���81�k# ��;�J���������]( , xcs���{�7�҈G8O���t+�y�XJ�#JK!;::Z|m�g{�73��!uO#��9Ȳ�Y#G��q�cfJ_���S��Z9i����N<����6�V�y�z��R����tW�{xl,�7�����kﻃ�j�6PA%�  �H��T� A	2� ���� ��J	CP��� q�9H@��4����}U��ڿ��ݭ}�nz���O��<�i��n��EO��P�,��R�|.�3�S�b5�@3��� ��-BvD,�8XPQ�Q���i5��S+k6��/�BUBpa�Ao(h�?b��_4��z}���E�w))�{�����sa�m��(�շ׀��q7��2A$�#���-+�At�w���-n2�1;>:����:�a��фk)8����!?wߑ�Cِ�b0ȹ\q&��yp�����d<c)ߗ�-w�{�J��Y,��<�ڪ:"D�Jޣ�OCK�qs"�pfNK�pesݜ�{�O���]�)JO����������%���WW����:��r��`Ik�����D��`�y��Q4u�[6�b�o�͝��s�2B���@�Q�z� w��s:O��t*�ݣ�L���祥���%�¶w�o�*o�������)2|��2��NL�Q�Me-X<�w^�mXXzb&-�9�N�N�#�*���Zr2[�I�dM��/ݥ�*%�>'i����dg��OK��!>�غ\���Z��kr������/���Cm�ӈ�Ly�����,|�z��!J
���w?>�}�i��eh�*y`�		k�]!�����4N{5j?���䐿<@b*�:E���BZԏ�w�4�����E/o�E@��Q����K��Kg����u���d�[?�+a�A�U�O%/���ϫȃ�E���Z%9@��o�h�l]�WJ�-����ܳ��*�yF�73�t_8�)�I+I�%���P���#˞���m#����\��_�
C�Q4���X��Ո�6�6? �@`q2S�a0l/�����O�I������H99��r���R�/\����c��w)�\��()-�6+y���
��/5ן���h�X�ӻrN���}R��Vh��T o��b�gdsgx>=��YK���dhhx�`������x��ƫ�v�f����mji�]�iV��`��U��	�PǤ��X����-[����Yl�/$�I�f��O�z�0�j佐���;����fVm�����T��8��뺻���c�K����Y�?O�3S���Y=�ɸ@��o9Q�u��4�dY[^�	��
�u��g�6��l=��\���\{#&�u�N/�/d`�}[T����9�[�%}�O^p�U�f����/Fg���r?~�,�|�M�3�S�~��*X��y�`��P�O넾{t�/�&ԡ��zzz�V������ܒ�7�����Z�շ���������7�|�۲��}���BU����[�A���y����*wIM�nر�4�ꈼEZWݶ�n		q^������}�M,mr�M�},�v"�js�!{+g����M��g����IZ���ƍ��8��"4M1��{����a11�ܔ�ܧ��M�b94�D.4�T%���r�,%��;r���AJ����o�q����Zr��6��&��A�����'����Z7��Np��g/)vc�\��O�ϑklGM����\9wGUUu��H@h�?�)�/�����x��7��T�&64c�^�F�q��P#V-V���gm*Ն�A8��B�l�S���n��������M���]���A��i 0"
8�]PMif]�ҾBe�GGN�'՝v�r�*E���6t�ϯ�ύ���9b���O�)E1��X���zs�p?{��t�lD[^�E�$)7�\�q�3��Xt�c�s�߈!](lcZ�b(nIk3E�^^���XY���ά������m�x�\v����9 �nB�L�D�6�p}�����WX�k��e���Q�y.Z������M�m[K�!G�X2R�UHS�Poxi�~���k3�/���55T�q�;����R��]�9[�4�9����*u�aT}�C�f�ze��]���@pp�bK�/�M�N�
���A�p�	ǩQW���?���0����8j.3�v����%L�Н
�&l�}��0Té�0^�0��KnW�6'>����'b$<����I���v7��.^��g\4����=�4�v�r�/�h�����
U���p�Iֱ�EqA��������RR���x|d���<3MU����n��𫦼�w�JdI��*oU�ĳׯ贋9S|j�3x�e��/0�D��=���fBz��p������h9'?����!	�ڒ'��H�����l���p ��#S��Y�s0:+Yj`rVI�|sCC��w�9杴�!k!Kfh���|�W��Ӈ����YS�q8���'c�Ԯ��D���ҟ��-ќބ��O��;��=_�6���wu\?<��'=���rG��ؼ)��O����N�1�嵗�0�*�e�,�L�v��(��|iY���년��./����&�2 �������!�[��/ڙ����b��Ue���h��b��$Qj�7���w�;�0.��#�Z�����+�h��7���?�9R��^_�h�A^�����p�1?�ZUU�<�r�������(�s��Yg�#ŉdWV�j�p��8b����3LY+~���p��3%L'/P�!�Dݫg��Y�Q�Wu88j=��
�B/���H ��A�B��J�!UC��0��34�$����������o�|����xx9ꚜ�A���@�O?��b�J%���nJp��������>B��%@,��+�]}��b��Z� ��Kz�wXA�:@� �Y�T��Cg?�ߩ�8]�pbz�Ò�;�_<F}�S��Ǩ���d����N�J���Uv��LM�{�z��ēf��~9�j�R+��|M��߾��ֶ�%��2ņ�䯟Rd0�ki���v��di1sf��݂?�\Y�Ys$��L��3�,�2�ï�d����G_v\ϟ	����gG��e_��r@;Rg�-�O�i�8�C	���������N5�팭W�����h��3����^�e�
!t��KnOU�����ξ�k;鵵�qO���{��V-��烊t�F�hAYP���837dJ[��S����W�#�=79����=*�UK�V�'$�y��*'�f��>�o�����(�d�������e���N�v��i��1������A��j �m�����Z�MV�
���}N���}����m�S�F����|i{YYY|��[^�S?N.��ә�$�9�,�?��s�4�qȒzx���4ɚ���A�ӳ�x2<y��wБ���[s(j��5���s��L�	j3>
Z�00iܘn6ÿ[�z��-�w��Ƕ�W�����C�x��)����j_���?�Ójc��7�%�	_��cC�?W��t}(|C~��"%>*"<|������緖e�Mןy��-r�l��5����v�e�q/�t�z��y�B���Y�ǩǪ�����j�x[�|��>��ܘ������/K��x�W�[�����b�H��,��_�d�ۗ�e�iD� ��킩�"�4k�[JA�wgx�����'�����ꄩTmLMa��o��'֚�(7@|(>j�~�]�����	 )ݶ�+�TW�ƅr��z��`�|ɨ�~t�Tο	�����۳����ljjj�7i�L=V�m�nd�cbB�L�����U/����_��Js�1�g�0���[��1����u"?Ǘ.��7�&C^O5�b�.:o�d��$[���"��iLLB�	���z�	��7~�w�����8�$0	U�zg�@��X_�Ǭ��T�*~�/�![�-���uz���E��n6XMr��Ϭ,��)����zC�|�"�oXr*Ϡh��Ή�ͽp�8�F�{'zztj�3�]~��θԂ��+�#�ON�}��������F���N���s~�x�{	ZMC;�w�[x#4�tI��M5uuk���� Pk�DNg���Д��P|�.�mc����f5���S��O��i�l�X+}(�|�"9�詩6$���|u����W�Y_��ؗǫ���9��$��"�O������_�$���Ă��N��O(w�*�]2��>T�'g�z����©�̀�+�Κ�~$HN�XM��MwMr�y�f�]W_��KJ�;����;e�+���wutz�y~��כ��>;/�arr2���ҘWT�vd�V�n���J?��M�����eS��Z��v�Bϯ\
�z�|�wB��ڹ�+��ܱ��;� ʭiA�y��Y�|a\�P�qhh'��T�忬��ʹ:�`Ɯ���l�� �jL�M?� kP��g�?5<�@3��sc~��|�̫!��5O�Z�̀Ȃ
ϊ�}��
S�cs�����dZ�@����;6F]�m����u\Z8�&��P���(*����Oi3�~�
W������rSsT��th����Ubݕ__}����K���R_���� +k��@�6�O ���3N�{ܧ�C̰�̑ryWY�<�ϝ`6��������@�o��j5�9��ԊV�J��&u�Nhk�&�_�/^@�5pq�%��3* �}|H�Y��&G���0;���W�㇤,�6}���n���1{�$�,#��B��o��U��禃�`_��|R�ʥ_ ��b�z�(bbcc�
������$ ��r��#�|��QPi_�R;�`�X9�Wv&�8���Q�ߢT?�$�%�1��>)r��e�UzEI���O55�}����oL�\�HG�<@'S��q�k�8T�Z]��q�0�R��UQq�ߓ�A�E�̂9?y��o�_���&�ȸ{���>�y��LU�Ж�HH��+�~>��
4��z��4���7 e����ʅq|�ˠ&	*�5<���y;sZ��\f����:�ӗK)ھ����b|�?ύ�4� �ڦ��7u㿢>7�������
��x.hJ�L^�"/..���$Oi3~�ڪ
���zxxX�QY���eIg���q!I�	K��%�"�)�t�U�AjЫ����ݳ����Q��	��ł���\�/:�t�T�ղ����o�Q��;�'&"�ހ��=iii0��Q֫ka�����m�ݫJ�b�^��+�/�6����[�B���q^�(# 9����u����`h��m�-�[Ё�P�,BI��G�=EE�?��f�,��.������?�n		Y�����%�[��
�Zu���J�֌iZ=3���kkz�+�M�g��Z�+�V����t�����p=/��nK��&m8���j���Ů��"u�u9���3>��-(��Zg�ߚ,��֪�����'���d������D����;wdd9���^�}�+�h<��.��������K�J�j��:��Pkq&s 
�Z[[鎪�7$9��t�]G\�~ۆ�E����kb�w�I�n���@��1��U؇��i'v�8a�����~;�Y
O_���P��x�~:h����"j=q�������_T4"��uVm��Nܻ���g�'}�@�.�[�P���1?��ʁ���Vqe�cB���>�b����(1�*���[����t�"�¨����nk��AW��?Ǘ>�y�K��w'�j��F�DR"�
��3�8r[ZR����ow�L9�&����6G'�ă�:�>raǇ�����r�3v�z�]�INW+(��N���	����?��:>���@*��df=�u�pHf�x��'@
�� :w�'o#�J\���>}�kkkˠ^�z���h�ׯ��P�M␉���ZJ3�o��O8����Bzx�����Gyo��r}��2�|z#CL�����X,�SM�]�k׸���1��CKO��J�J�i壽�c�5�1��Ǐ�-#cJҘ��Qu�3ͩ Y�轻>ߡ�mO�N��l�BG%]om�F$g���Ԣ�,O�w�K���ߐ߆i�Dt���:ZH-�l�&�G���Z����z��>/ �@o� ��WMߘf��+��Ϸx������!����jo��.1<����|8���������������F����?�ܿ��rʷ��9>������.���`�c����K7U��Z�ݜ�_p7�:Y�x�XO�$\�-��M��jA<n`:��/ak��yΞ=��a�{!�Q\R����X��s���h1h4z/�x7ꀄ=��'-����:��Jv�C}�{�<B��G���
��!!�x՜�g�"�=S�'�L��/�d-����8d�fƽ&p��{�5�ۣ	h��bꀃx�ׯ�@���rq����I𬶖��N�[_���ǭ�:zzzWW�7���''��;Mt6s�')L�I�K����MTG��W�4�3-���pmm����cv�m׃�m�q�)����Ԩ❍T�u�OuH�M+��z �<'��%	�&�7<�̮�
��r�iE�����㠣f���'	Z4��b|$�Ǉk�@���1>�e";QC"�t��a�k}��^Q�Μ]b��|ŧ��Δ�>�;�ܴ���5W�fw��2���K�5︮�RJ�;p�l����V��ks��}U�'�z���8�x�Ǳ�\ve)�N�h[q���OV%���:����L�i0߅��]���544\fg?�r�U��G�t��M��Z�&NV�qK	�P�(� �BKS���Q ��o#?�\��U�m*+J�u���c��%p�K��K�92'�晰���(�
d@�
U��k�j��;��45��F4=����&���2�;8 ST?�:�<Wx�."" �+�����J����`���Byi8��Gy�}��}���*�*�7��*��̬*v�y��4jb�LZ�����ph��9���ŕK�� �����<.Зz_Q�rz���꽃�.7 �yLT�u�C���$�}l�Fᩢr4����r�P�d
���t�����ڳ���pv������Ǝ�CL�_�o��׊,(wo�?�J���#��G'n�l�v��_��t��Zk�JE%��#�P�Y��2�-��A�AN/���|Y�Y����12�F~1��ӫ]��ӫG�*�^��7�J=�ӵ$\��#�':֏P��܀n�p�\ZZ241��L��O�,��L ��C\�]���SVnni��/{�d	�^�[�a/.���2Ԗb+�Gd妎���5�؉r�"Xq�0���a�rs��WI}>�Щ�0�6c�;s}�!V	�@����Y`"�vV�ۓe�\�����~R��������/(��`�}̨���>��7�L������ĉ&����.-��Bd��w��n`����+	\��`���+���A�����VSs��Is��� <�spP������ƒl/��l�z�j�uFd�;dn��ɸL��&��g/��ɶ8i���<1�ٚ~X�P{Qb�KD{�m0IU���S�R�~�UU�D"�pW�ã�J%_''{}|dXYY_ .^�����Z���4��\�s)̐A��,a�d%o�n���Ӂ�kTP��
e!L����M1
+�_ëZ�H���z��j�|H���t����a�wَ鈣Z���4F?O�Y2`�'ة�2|��7m�#j����M��g �Ŷp�ט���!�b��/���\^��,*t��	\*b@���鈝H��=+n����s;1��<;;"5�,�*h�lV5���=���LLǿo(0(�_{B�555��r<d�<����Y�6���I��Y���4bn��-c'�ȳSr�[�U���l�&,�a�1�vz�E���=��KIIĘ4�:�s��PS{`��Vh�^�M/PT�i���4���!4("�c���9�K�ƖjRjJ�0�����S�MX��f��?Z�](�j��*���z�sI0VC�yBȐB��'���������V/���zP=��;�堯�V�:g��7[�v8� ��^���V�ě~(h8ԠD'�ʵͬ_/i�ٗ�#,��k*}pT�����W�^�H���;e�G@���3!��[׭�*Ѣ���zzz �o'���Q�Us_
����kC"�� fZc�0��Oh��&o/�[c>���V��o���qݝ�ie�\@%�ɪ��}��9W�.����w��)I$��x��1�I�+u��\�����n�� �-A��{ˇ�?�0a�f,�uR0ǃ���Ta���-I&x�������[�ܟY�X
� E=L ���*���}�.�]� ���R/����~�٦ �Xa\a������$�n"<��їf�(3V"Vz���GC�{��rMlE��+Pi{�G#����f�uia��rԩ������^㕌�}W�[�d������'n�qs�$x�v��hf
�z�<-@�/w\
�1v9��=h�eg�=�F��,#8��J��4�x��v��k����P?�i0�2����ና]�D���Y�"�/�C�H)g��j���+=9���x���,<��4����,�� ;oU��t�`���m���`��ziZS�= �?��U�s�A�=��������L~�O�n@�(���l����cd�\���5U�˂�d���S֏�/�L����.�@���K�o���L�#�5�/���4�p�t�3ܦEk�8V�g����VC���|`���y�J2�*YS��&R�Ԟ�D�S�`u3���"��Z��m0�W=��mbc�z�X`�&��shel2��ļß����s2�5}�36�1����.��e|����ϳ��x,�Nn�f[��f��u6a���յ��R����`��88@�� pK�݅+ ���;��4��Vp����'`�Q����$փ%a��:D�$/��.)�d���nEn0�[%<o�.ic�\Ztˢ�z�p�(���h&E==���'y����a�A�Vrɬ�c���I�t� j	ʄa�XN.n��ڻ�ᩃ�0k���tUet5��0s
�m��b��MG�[N"�As�ڳ.*�6���NDl�w:_�w�y�]p̄i�7��P׃�f�Z�ؒ��f�إ��]Oӕ����G�����f,���+��&��sEH���ZEmc��R-3���X�^n?����OZ��Hl��?�8����e���m�L����e,Y�������eX]��i�n�n�p�71�C�}8�>�|��N˯���\iL�i ��4�䟼��G�U%�t�"x�6��{st�G]'��'�������u�1�`��@�p-��U99�SxD��{I(=������S$���`^��	�W_�1ǀ��F��-���f&��$T������}��Y�TJ����m�9�T'Z��9B�0}8�����e�����-�����W�S�yHqT/O؎h,u�i���h<���1֣�rM-�M��x'�g䰮7Z��:7�#�\s1���vE�W�����ǈ��	��	��;g���p%Fg�dD��X�u�� <�����1¾���M��!ĕML)a�� ��� āh�H}h�@d�ȋ�s���o�]>=;̜퓵�$���P�aB�늌qs]�mx8Ǵ�Ͼ^�<�g�P��,��7}���x�CK��_������)�6����~��$t�MB�3}�m������;~�	��|\��Y��ȏ�9vO�p���+d����ui�;�`�mґ�tDu����[$#l>c��^ʫ%��t'������8w��i[�t�HT^N����\�28J�����\=?|��fM
���>�Im ?�'�g��ȧ���z_��֓���(�Ubw_�U�5�^n���ʡL+�N�]i",E��NrVP�������k~V�`�D'����l��=w��gݜM��.��vy�X݉��(-+r��>���l���->���g��W�:?�i��a�k!0�}��Ʉڙscd�v���o����&�H�0F,�ٗ,�ǁ�����K;�40cZi��}0C�550���2MT�5�L���������o��C����Z�Y2�h����~�ۿ����ټ��9n*�5'�@���׼W�d�? PK   �m\XvO�XM�  Ի  /   images/6bcbb164-c8eb-42ac-bbc5-5fd68c68ea6c.png��S��=LHA��eq'�%������!�5�[,��.\��	��%���_x~{�jj���L�۷�t���� ����g	T�g)�^>=�/z��t���ꄂ����|�ȊC���,-Vs��o��B]���Bu�+<���ǹ�c������%���E���?$4���['J�W��]7Ë�3bq6M>��7��`�њB���*sO���b����炗=Q�ȁ����s��ǽ�ɩU�ͩ��T[^
�Q�+�o����4�R���Ď�׿�W����I����0d��]_$�s�h\��@����UK�_7.���)^l���W.����Dh([���8�<����kn'�������������K�)��|K�pZ�3I�m:i���E�䩩���Yh�| �<E�4E�7N�9��0��l�gng�2��6Z�z��D&i�A�TQ�R�3j��\o�-U���@���.�e`�!I�z�j�V*�Á#�[>��B�J�k���+r�e��x�.�2���i�V�� [�w�,�i�6��{_�G���M�fruq���N$�ɦ�B�r����{�}������/>��W�o,��㹡�������'r��Ƀ�^X�]��T�]*6�����r���+��ʙ5�9���n�jҊL⯻�N*��j�-�:!�#� �=�gO�Eʡ��V��]�,�o�F�ڹ��z::�@���L��r%_W�UB%	�^�I��i2��CT �I0�lܩ�y�;�O���ѽ�u���zr�&?�Yg���LJPKx/�IP���ߛ8�F�!o�Yh_z�/V+.7x��i�y"�+{4���.{@�ÿ��;��P�����gC$vn�g5�To)(��ڢ'ssseJ\̮޿�.1vMw�2�l���˳R;W�Y��~��Y\�h�����V]vP���Y�O�q�kQ?�Ҹ;Azo�
t�V�6t�,\s�S�N\��O�5c���yʼ�"ܛ?�Ve��R�؊����ؽn�E�v�� {G�o��lk �ZD-,"rG�)6H��������0kKKkR�,�����s��kۦ��^���7ͅ3ss� O�Ȝ�y���Y�<����\���0�c�����L����|�_�	쨒�1E�������_���N�]�A��ӽ��:K|�Ͱ#�����<�B��+�����d��k�co��)w��'l����f���~������"&+t��o���c{V�.���G�&�u�����g5���K�1���b�>����Pb	z�/�_�_\�-��{��	���ֵ����K�������p20I��:"�i{�y0e�i��n��e����Y��:xΣ^'E�=�*��/�(�(T1�̋��YeL�ރ0QPjXx���VL_T}zݤ_��ET��:��NO<Fwl00��iHt����}�r�����D�Qډ�l�	�4Y<�rq'�q�]͏�Ȫ|#\��1e[?��[||��Y+��O���V��@4�*h�Ěb��ǅ!�h��Ӓ��NjE�1��,u_;5C�s]^�5p-Z���t�;���V�x@���/\<כ�x����K�;�w�߯2f�z/"�M��r����)X@�+*��#��W�m
s���P�eS��8=�nC�{���i�t��a�p�'�*���1/�x�������o#w�sV��֩�����ۋ$kyd��F�|[\���@�G�eoݾ�����z6���ٲbU����H�Y���Ƕ(��DC�Ԏ"���B{c��_��K��z������*�U\�"F���M��p��* ���XH���^��޷X���'kD:,���1�i��U���e�A(����;�)�����c7��Q�0^�S�c��}^��FmVJ��l��n�$�n�x�;�&빷*z,�_1�9+uU���q��xB�䮋1e]Waӑ�ز�@�F�Ć���
�4;n�"x��C�.Pz!���u�^� ^lD;2���

��21����'p%M��s/w<�d3���f�����M>²�s�#|G�c\�g�M���j�r������-�@o�jup�z�_�UX[{Tu,yk"I�˸�5}]����J�.���V.v_�M�8��U��2a(4���s��g7 ־<���܉���S�^2q���|�]l���1$g�;�NS��!�A�cD�ׁ� R�zV��}=̠�����|�q�x��	ZeR3f��������Ud=N���_�ܝ�Ju�3��X���đ�h����ڝ�#��xڙEm����ASK� �ź����}�濥oʻ��G���"��'o��x<0�K��H�ޘYh�[̝���ὲxi;�3ۛ&�K��ҿR@�E#+I	�Z���`�B���S1N��I�㓹<�a=8W�O!_�����`$V��r��d�	�O�������0Qf#p�c�ڛ� Y ���@r����5�^")���7d)Z/E��>f�C����~)�,h!!v��'��p�߼-(�֗k�1z*Poj���]��z0�ΐ�@�(z�O��M�$� h���-���Ը�(��\p\w7&�V�].����_�O�
K0�4�=�Z���r�g�+T؄���Gu�xp�:��^P��Q�Ą_��t�@�#�l#��&.]��qVJ+����e��Bz��=����;����9nȵ��+E�%������.�����_��Y�o&�m��İ����S�ͼW5͇b�r����roJJ�5dh�iN�VJ�`a�X(=~q5Uzq>XU�	�a���D�pdp�Xè7H��w��5D��ʩ����O��5�'�DD|��1��jI{���j�p��y`Ǩ�;w�!I��Y��м.�k	Ҝ�ߢ'��ý�����&ˊ��?w-D�'��������X� 	X!v1��"�n3�(�f�����g��1�l,mKe8���K;F']&�La���:"S_E����TSv�@��6�PE�%�����m���}*�#���RZ�&iC�'k�ff�����F�%�O��r7�,��na��f��5� i��t����;��'�W:�X��w���'J/�t��e��Z{k.���F����N��r�G�5:me��4�V�#O��CN�a����׺S��`�WO�My2l�6U�:T=yܒ�����ĕ����!K���z��V�7�k2^�-vt��-4|�����Eg�>J��$2����/��KW�Zb��@�����C�]����Ϋ<h+�j�B����ɮ���l~/�F��~K���4d�'���o笯!$Ύ���|J�+á��9zL���(��%`�|��f�[Ƨ�!))=�����^k��ym���Ǘ�`2�֋ԑiS]�mG��L�j�-zZ9f� "plP��N4��:3�w������L#�����3�ܞ�bV�����}�2~�Z�Ȼ�P�&��|�/�œMg`���x+x��e�ڱ��̯�D}�?؎d3�rO� ����	nV< ����q��^��y�� ^} ����?Ǥ����Me�Dѣ�I��UY�=���a��)>�.��Ljܐ0uۇm(Nv���l���d\j���krc����h3�[-{a_����mD�����hTUZ�6�׭=j,�UW.D8��u.hWܡ5�r���I��℉�����0�g%��F�Q��#v��~_*��ϡ�ԧR_�jӊF�oE$Go+�;.���lA��ij�,�MmqW�d�X��CYo�rٌ�Tm_��i��_*����ҡ��)4����]���l�������v�D`Fّ"���}^�ܯZ��o�⣷��b2*�52H���bhŨU�m�d�	��K�P���6�4��aٜگ�X��b���M	�	��������Xc��/|�`�F�v?0��ݓ��0�U<)�O�]<�Q�"����h����Мou}�s�����S�^9?����{�]\�$��/���Dτ����=Sl�?;v຿'�Uc��Ң	|ù[*<Vq�2���U�n�5�Ԓ9`��Ӥ�Q�S�"��5����q��-�$.5���i>��g(��L0��6��f=Nc���߮唗�� ����q�:������Y	^Ĭ�E��%h�H`����W;�iBe�dB2�֑�4���g�@,��SML��!�F��a��A���<a�@�W��[=_pȱv��]2Ў�Jͬ'Lk��^Y�;<����j9��q[č"�'P�sm�97�d	{�,�6�>�~��x���U�률?����v0�J!L+�B�BB3VՊ�=d���&N�/	!�|�/�cI�ۀܩ��\)]����
@�#����<g��v�U�Y��)��bHԋ�AW�0L����v�)wN���bI���'�e��HIm�pQи�||s3���ѹ��َ�����f� �79]��M���0�k��6��(�����^��z��͈���٪�=^��{���M,�}��Y+!l�F׀!�d���IR��L�������������mv��Q�wH^m�������<!/�,�Ɋ�d(��#>�18�����6����:h��/���s������R�1� 44d���Եut_L�����>�8�����V9��hiTYfV����C	�;1��^) ���7������S�u�\Ӯ}�s�9�Mޞ��^����2����ʩݲ�&&�ti�w�ّ�N콶�yq,�F��Tz�+dM	�I�$Ǭ�R�s�$�������@���5��>�欍+�d�����
vaAa����1�\��.�)+�Za���j�K���7���B�����]��j�j�63����Wt�Z{=5����t�Nx\V����Ol������l�/p��1�:��"闧�a5oܠM�0�ۄƺ���W�[c����G�E����:Y�;��KF�0���&�o�*��ՙv�}_3S���z�>��&���qhȼ��GmVi�eփv�a�{�b��	�7D�ui�r�g���E���h�[�������枏�'�	;���v'��f�8{F��'0�&ݢQS�����|M[�|�03%e�RZ(�lٶ#//�4?4�؁���W*�j@0���.�T@�Ħ���ZXz���$�H�H�bv����~��J~R&���U3�tי��2&��M��{�J��(̝���e�lm{k��� �\�O�#���>���6���q��R7��5TB��6EPP�>��Z1�jD�uv��Y�����F��RPd��YDC�ݶ�u
Q=�NaP�a�L�xG�\���i6Vm��/����t<�jFl_{��j1 �=�����7'�������������?�ث+��<�Է'54,L��E+yߟ�Hn�$sl��M�5h�+�&Q0�+-𹵱���l�8�$��*���B���Ő�a�tלq+�k�݌��Y<��q2�����e®Y�����X�7�D��$��f%���9@�gb��g�v 8��1,d��y7S�s'B�&<�Z�l�����wbC��DM%�����ykk�8��&�"���A�LFӴ�����+����a���q�QLDt��h���R1>���z�+�k��w�X��*SWӐ�1<*=�c3,z!��E�8y�4f�*�M�#�ܟ5�e���fe����w�Lo'j��+d'�[������t�F�oL2��cx�|;.~���������l c=���n��f�.�͒6��2��t�au�����8L����ʐS� %��@3;f�_���Q������Oq?����l|5��`���<b������3}m��+�����'�a�N�z37ޯdu��m���ܧ�k�m��������@�)l�oyˮ^[�+w�K�����7��&��N�Ek�����U���?�e���ڙN���Ύ{��C���v��[��%��IeW�!����E�'&����3tZJ�F:֟����?-"��Hq$`Nd}	ꗣ�,�����j�m��d���*dF8��UM�|�`@�����HBWҫT$��P䫩�D?�cɪ�ݢP��FZfܾ�F�I�����\g�� q����)����S|����I��BXc����T�����h�쯖r��$`�^�e~�獷�����2����p��=X�����{=�=��3�­(���C�r���.�����7u��j>O��o)T9�é�]xb�Nk���>���L��X���[��[�$x�6����,��)%��$l<o?��t��}��v����o�y���´��Ҩ��X���9-M9�u��kc�%K�d�-�@���݌<�
��<
�x���A�qH9QZ��--U�' ,���S���5�]ͅL[�Ck�tTP<ƣ���/�Mh�眳B�;�W�V�H ��'�AU��c���'�;����s5�����[��㉎LIlļ�bC')�ֵ��SVf#\�%]3��I��l��8=�� %�1�w)����������'UZﲀ��o/o��/��(��Ǘ{{]_��\��	�ͮ�q{D���Lo���Ê�Ϭ`l�{�g#@��a��n��?��D��7S�M�䟂[�a��u@7&O�S�X��-�4D��ZOiy:
���C]�V��B�֢M���@c�Iգ���&��E�e:�M�TN�8Ǥ�fױJ\8���	���[?,,�V#��'s��O0��o��on�Ȏs�o����D�Ld{I���B��e�v<\�R�����ʹ�d��l=e��j���Xp~�$M�w9�T������=�݅$6RN(]	���G&�E[r�=b���+.8�fj��h�c��L}2E���ן 2�2���5s
�F`o��Tk@�+��6�'8�"k"��e�;�l�0Oݎ9E���A���7���
�CG����F
a$�9�0��Ll�� ҳ��,dh�F���=X|��@���1�#5��fb�ޣ��i �_c5tQ��_T�����@��)	:����Is��`z� �j�gxe�3�aS�������1��ZWqO��t���A���a��⦙���
Ą�_��:�M��$�P�M�	�p�^ו9w�ܖ����:B�[�y�Ob?�P�����<6��_l��d_��zoj=�WX;67��(�h(��͘Xx�:��7���+;�ė���Jw��	8�6���~��9�����n�"�h��4{�o�?��#�u��t����� ��[]z:���`�V_���a!�I�nM����W�Q�Nh�9���?mN�$�ׂ�P�����������h�t 5�P��=�V�'��F�v_ �(�����CñϽ��;���f�&�2�k���`���y�4�;I|_(2�'X����^22�]Z6/�|�:qX^Į����G���h��c-XRg隤�c/�:�����0"�"_�Z(����%Jr_�*������L�֮y�}�/��� ����sT�IO!��Ĭ$�������eR�GW��X�6ES�}�@�C������zi��� H&�C�y<Є�R�أ���;2h!�o��. ��w|�2��*e[r({E�}�+3�gwM�y��Z�P[��i+����Zls�"}�p˜5��pk��-�RC!*�|�z��Нt�%�>{���S��#�MQ�v��:���{ykc��_��ō��anE�NX��s o$��vA�ֻ�Y1��t��"�8s���SCv��N!�gDHĒ�)t��E-����L�,�龉���ndD�Fi#�N��z�n�"9�aW��_QV3�>�v"e�^R��Ԫ�[nᑂ�/{X�����Z_����t����-$E��l��3�f�W	�m��e]��m�n��ƭ0RљR��G#Me
��O;|�r�MN�Hw��wl}��"n�x�8�ˑ����:5�ޓ*}���*���:+�y%�^�F����zOt�u���e�tl|j�'�P��=h?�Tc�"4��Ԅ������moݠ
,��=�n��	D
>fP7��Si0�	&����8��O!�#��0Q�Y��a����b�,;/�['���͜;�Kz�G�z�_��s�f��ףp�\�wv%r�?M����ց��_&F�z�D^�h�����c�S��&�Xq�ʦ�aK"�g�-�,3�ںZu��3�
+�m�?��Hڱ�����r���G�a(�}[�Aa�~�h��bt0J=�M�gI��_Sέ���V.qj4�Ό�[;6AG1V�VuF!��e��@̠����P�p�.w��v��N��^��\%&��<9������k�6�N���{g�t���=�4�6W��}OO���@��]�z�SB}�٤6�T�Ti�_��$i�����tXmR)���;�'1U*sC����/�c�mE�z�*y�M|1��]+Qt(��T�.��P�NB��=�n����l�z{��h@I+h��<�\��ښU ��J��3�Y?&M��{�"�D6����c\�`��h-����П���	�2<ݽ֊
����D�:: ��L})�r9*G��Z�8����ڠ� ���>�Ghh<�2$}��d�&��(�����}�w�k�)I���B�:1�eQ#O� _67���p�A����
�dz��$À��W�i�iƆ���<�Ѽ;�wJv�}� ��Gj]�Fi���za�ǝ8�h�X�:��U�S��(hC�wY�aaU2q�v�*ޖ�s[M�/I]m��,ϲ���y��N7wp���걠��o����������{K����_�$F�&f�瓍���(��.��k[1wi%u�xF�U���,�=\���ܣ[�i����w�㌊�w�{Tw� cŝO�A�[���f�@\H�Uy�5Y���i��/�T�[�!�YXtV|�c�$�p����j��䌣9f��^=�Q��:�ztM�H���/�K��������y���hWW��V�?�OG�遽�Wv�8W��Q5�*�5n�&b����������3?|%O���~7��/O���_{'�)�	
0>C�@��� n�J+N��<c/�L�(�N��N���rQ	��o���~��K׬~��ѫ��ⲫ���Ld�ޯ�:��V-��D݄���f'B�C� 規��A�����و�@�Ar�q�N��͙Ru��!V�G�� ��(����~�摒�Պ�g{w�|�Y�/}2��j�~�\��( �q][���oe�o��W�n�N��o����u�\QZIl(��=$M��ۅ(��v����({8Ȝ�GL���R!�f�A���j�z�U
Ly�Ҏ�w��ҋ�~��b�7���(�a����u���6�.���̏,�O.P����w���[�_򶛊�9��٥�G���w��E�D���� s"i�ndw tp�vn���.��qM �m�OD�,5'9���/u�ӒwT�_�g�����\!�O�s���q�En�Y'-�o������q�<
�3�<��'��>*<�K�-U�Y��B��m]�����?|�Q*"�,i�x]�v{�.)�a1�ki6�����W��>��0.G|ݴ��Wt]B�e��spl`��-lg`L��EO�c4�k+<[Yn�
[�;�d߻m��z쥺˭mi1��jm�i;ޤZj0���/}�̋��%�_�wv/vF�z��t�D�W�����H�c� ��kt�����N�V�.��&�K�Nc�r���-1�E��yI�7<g]��`�Uu��E�ZѺRU�(���-���1y�Ma��bL��J/�v�N�ʌ�C�{��Q
Ә1)W��,�X�v -n=�a����[Z�F���:N犚{Tg'�ae�̷Z�o����5N��E�]&5�X&_*җ*5IL������v�1A���O캷"�%<[���������[��Ŋ�B!��G������Tm�/[�O=�C���9p��)G}�f�i�%�ȇ{�-��ݻ���x�"�G��V*�H|��\�6Qo�W�Y��S2�)�g54�����k���Fubs��(*
��������Pݑ��R�r�x�xYn|�9���[w�Z���\���K1\��%�ӡz��T�o�׆� �N��پ�8��[
}Db����%��o|�D^û��[��d�n搤_{�Y�ҩK����g�J[��)���8C�G�(1���z"��5�(�J�n�:����s��	����_� �כ�э�Km��/�~~~{+�����J%ZTj9�������g��Y�_���c,�	�����s}��D��JVt���!�=bTTk������,�2.�v�)���Oz:�SҾ�A�Iw����z΋�,���5�6*�#������#������ˋ�>���Ӿ��k~���E�����{��[\\���{��O��wFE��nvA�z����mT���d�NYO^r�����~�U<�Z��'��t����7��]W���L�xy��|~V���O�l�zᦑ�#eTI<di����Jg�3{%}&u((��E��n��� z^�lŐ�Dׂ�?����^̞n�X��6=�D���U�nn2PRP4����go,���i�f{�������ā�kqIl"�(Wt�a�3����RO��j9��I��4�U&irU{ך���D���"��q$My��I�WOJ�i�[��٫'n����m��=X���蹴�[���X{Xي�����*��"FOY��=����q�$M�s+�46��ZK�<)��L7�hj�(�J~,�7VqKd�e����II����fy^6�x
I1�N��Kym-����ʹ���<U ޻((� c��c����=�F���޽�y��:���P����ߍ�Ø���0���|����\�xG{a�RK�ڳ�+�Z����������S�Я�̠Z��>D�D�k陝7�C���0S�|���*w_�L9�%Q��Ŝ53AJ2j����æ��_�1=̇�_>g�b�9�58�[��fP�Zۺ��s���:�B��͵_�]]9:��Q�NI��j�矈Ѡ���'J�s�>cB��.�0T���֌�t��?ޱ��d�ϰ��98Y�e�lY��,�;X#V������pN�N/�}�2�DU=DAz����`�G�ȋ(T�E�+�U�|L}���(������I�L���/�>��"<C���Q��μ�2�� �c�'s������k�CX���5*п?A�>� <��>����ߍ�
=�G�kU����' ���	dZ��껚���R��K�Kww���x�� 4��/d��eJ�p�}U�I��P��o������nv,�ZF��Q�>m�`�)B+�Yt�*����TY��^��n}x���O��̛%��,��(�v���momYZ0���q��T�ǻ�]#fjU���n5�&�U�O:Q��v���v�f��ux�M���ּO^[ O�R`
�q{#���I}��Dk� s2V�XlM�p+"��o_��SO[�v<^����郍;�����t���P�3hhc1��K T�LM� ������`�Pi�1be����4�I�Ӏ}�yI5����H�槡%��u\��R<%(X�,e��+!��Ћ�0ZENK���x�bPš|��h.bVFF�v�~%������_Og����a�@^��zi�J%�L��i�o9�ت?$���/1��̈́%�r���ib�T�7�V���K����f�wFÌ��dH)̜'����T%#�>4
YN��{��55>Gs�D8����W���
�s_5�a�**e��2�Z��{%���O���wz��ͨ��;Q X�ˍ�Ә�%��.� ����R+I�d�|��12���V��L��ОV���H����T4c�k��NjY`r
q�Su�cB�<[ۤ���1J��~���`�ڊb�H��xj�Y��np��}w>�w�ܓ�(���s%��fD�`��V��}mQ�J"�xR�+�k��U=L�E���l�_�엢��n�Ew��r��⯽��	Â�skV�m'��N�dT���6�jC+�K:�A�gFW�(2��$m����&F�ѽ5<�i!U�<�{�f���W�Cڗ�e5��0��T�N�j��66���(���t͖6�@ ��������.s{u�Hx�L�8�F��+��JB��GGg�����p-�P�;���ǲ��nr]�O���V���C������#'}Q3�&�{��喥<�2i��:�ߵ>���eݜ�5���y~jٺ��i/ܻ[��Gr�T��*�8�	ns���M��G��_�k�
B/�b���;�Բ������kR����*C�a�����턐p��$�/���n�ۡM���s7d��.鬃Z#]���4u�|B��G����ƝOݳV]���ǌ�������k�;�Tbo�kJ��2��*���]��R�ߛ�B��6��r4p������ :K�M�����	��R}������?iU�9�%��ԛA��z����r�Rv̢�aa�ꋁ�t��;͓G�ż�h�Gn��w�='3�o�nZ�3_�LY't7��i�*�@,a�5կ$_ID��g���M$[`z��'���*se0��4����~��А(��M:�:�Ľ!tztf�|n<C�r��d�J�8@y~���Y�FL���*=��v�)��PM��_�D?�$��H������;zz�������Ֆ-�w0#�ѱ~ɡA�M����¿m*�ﭯwi���'~��	
�	�*�%��$»*�?K��-(`��h�J˹Ig�<�U�oD��8ϛ�z�+�4� ��1g!�g�~���H�Y�F�ݘK��,��p�֯�*��{�k�%ٖ�gW|���%\� �w��^�3��Z�4f��꧂�]��5�Hm�N�j�'S��ǂ�'�(ur1�k<��&�6���d�
��Ĉ�PVNXT�E���T�u+оi��X�lv���:0�:+�p��n��c�4m��~cv �ִ�t�����!u�6��}�+q	7�m%iiQB��3=oG�H��p��ܞaax�F�ݤ�k^�V���k`g��:Uz�iJbx�DQ��̵�D%�?����(��&L>4��&�*|4Ts�w�]P9&��9d��1I��^�UWmh%�'���>H�]���n�>3+K��xaE�1�l����vw�e~͵��Y�d}��'~�|Q��[?k UFK�^��M>���o�.�<�H���W*��=PA�o ���Vڮ��I��H�;p��*�ܙ%b�=�a��z���T��=r�w���K�$=�_ޛ7�֮�F@�LpP�f�� �$D�y�e���q��V�+0��-�!�KG)�VK%84H%�x�������_6�����]�:�%*J�*������=�+���j���βC�l�N`��-�������Ό84��Ӧ�F�*R06AE�"Ǧ�{1@��['\�H������^�:�7�+~��;�X>����>>>V���/�D�"-�t4���6�_��s�����7��7Ś�]ϧ��\�7������r:}�?Ҵ�
[�NM�܊��Z�M���{�N�yf��v潇1^� ��@��:w)q��((�L�u�+��f��k|��F���j6A#Γ8)���6p(f�;`�ַG�&M�p���90 ȏ�4X�(3����B������3
��,o��-�1��N?��UJ�G�Uw����Y:�#�p��|M�^�Ve�v`�X+���kĞG`Π�.����X�������F����T�u�rtwgeE���T��U�k$k�.��Ӯ�c-8>Τf!���%9)�l�gy��6�
_��ʬ����9wVK������*�((���7������®����܊:W#'U�MT�M~�T:����3�Ҕ���.�w�yz�d�Y�BW+�*�JM9���9�YS�އ�EP7�w!8\��X �o֜aXV����/-�E�U��b���N�U��bF~�u��������Q��>>�U`�շ*U��3��{~�k�h����j|E$=Z����p�b~�[��p@ā��F�7�7Rb���p�"�%(��[����{��tD�\\4�db˦U��"�ؗg�G�q��`�*��7�ĵ��j��fmp���7Ĝ�r�]G��h�.��>=*�,���W��Y,>��TU��Qv=���:��%o�su��1M�{n<ߦ����oJ����޷��8B�8��{����FN��Į����|4Z�o:O�����Y����g#�QQ���>57�ɖ���Ï77#V�H߫ 1إ�IV�����ăs4W����|����K@�L�*= <ֶ�ݑ{U��������~]w���L*�u�0E�wAg*�v���ſ4pJ!!�
�:5>�,����L��q�ĥ+���!��b���!؞�`��-��ԙd��+���4�c�z��_�vK�H�ծz�~�$*���r܍���2�V2!�b���b*B���-��YRm>%����վ�;�l���/ې�����ϙ����9�_xWƺ���7ec�������&"��.�����Sy�hLg ���te��Y)�lPM���`i.��ƕmp���X ��$f���|w��i�0�De[��k��)�v���P5��r�rο�����g��̘�Yb���6ʲ��,���O&&U�ʁ(=�Y�����b��~��;����-r��)'գ�����(u��p��p����!�hZ���[Py	����!*½��~(�֦�� j�:z=%VD9�� H�B��Ƀ?9u��A�a	��� �.���'��>c�8 ;6���� ���^Q��W��h
vJ1K�|�	"^�'��'���h͙����4�3陭�_ ��AD�T1dd��:�C�:��vw`���[�QɈOGh�ш��jN��j��8�������q��}sQQ4�X��Y��BUl&��4b?����"&T^��"�L�A$�y<���ʵ��=:YP��y���~�s����
�WUK<�p���e�ǸF��Zm_w`(K����(�md�-�Їe֓�L�2:�v� 9��+�qR���p �Lk��5�>��tޓVf0���R'2�{�B}5�G�Z�wV��MC儢�%'��DI�y�0�-�2�Ai}	o6��;�Qƭ74f��,鵞]9fb����^���(���c<��U�w�,�<�-�������N�E3��d�1��;��`��"���j��,���ױ�b�����-8���%�@��6�A�"6�).<�)�$�߶�1����OEm���Fl����v�y���V�q��Kg�勇��u?a��j�~�w�5�9@�:��a�c\U����͖N,��$���F�VW�7�dY�J��܇�һֱf�/�<oi�h�5#�����a��M��v)�)�a]4���RB�l}E*�7��>�W�4t�{xb������υ��˄�iҷ�m�Ya�1�b)�m�tU�vaL���<$���_���1��"�g¹f5��Ő�d�T���FTi���*��x��$̊�4��-`Zu&�Ø\�S�W-�5!V�5>)�Y�'�VL}fV<dA烘���}w:=�N���������A����7:I(_Ѻ�p�fP�N�:�b�L��j18N)�����'���&bqo�&����.����ap~�
�1!�d���������El�ƺ�7D}�Mw��WO��x��ª�uҢ�(`q����I��~�\���+�����q���Sh}�9Ia	��6,�h&!���S�qt�c��H���?T
?@_PXHo�&��[�'@��Þ�����Alr�t��Gpi7����ZP����NIùo��m�7绁z%��q�H�wg#Qx�9�[@�x	�̓�@U��4B���mO�ӯ���0�ı!�qu%�9���V=�4��̂-�?o\��4ݐ1��U�%�;���z�CAx^�\L��V��Ag�j�v$}(��Q�/��)���:�M�57�� /#](�St�)5b���]�|4�Z�c{����͑J4^���#1 �����x�EEz��s�a 01��#����.��mN�(@�cØ��0f�.1�Y?R�����ɬKcP"vC���Mƨ�R�N���慥��/m��>��j.���W�˙[eaN�agN���რzG��62�[�e�~.�����y]p㶘�k���@
�'7�@����D<}�ݨf���F��鏜��K-u���z�Tˌ��u�U��T�����gڟ6K+�����!�.�_#C.~I�Gϡ5���j�#H��H+׹�ԙ{!}�!�0q��c�(�E�f>�&�"H��Rv���&��G��S�/|�.Y~B�>���zn/��ZWW����� uy��X����~'���J�E��e��$����Y�Q�4��*����X�Q�2c�=��^��E�g��#�*�궨 JIwI��� - �ݝC*��P�"����������'�^{����sH1���G�~�@{���9�4�C���A����ȥa��?�&�$=��*�\,9������ma�=,��/	Z�ƞ=��iZ�xM�7�Y�ڪ�)���1�Qg���`�Fa������ë��1�����aVh�j���G|��vƑݿPc=�~D�rj�D��ց�/:/[:72BtUG�wWDM3ޞH�i��4�@�\^����O�!�$�H��NZ�1a[8b����E�MI�g������o<�E��j�V�Xۏ7߰� ��5^�Ӱ�z���1�A�lOG�I|��x�9 �q,�7���7�YJoG�\�Zrb�r~[Г��Hܰ����t���eX	���CC�:^(�AeӋb[��G͑܈�ŀ���2�.�;��o��M��Z�爩e�i#Zce���l����/�^�\�[,���w����OuʹV
1#����Vӄ��go}ԧ���*�46��ȤO@���m�	K;T)�DDD'''ϟ��W����/N{Ènu$�6Ze`���5N`�m���.+s�W���$�f��A��c��K�eh��7?��`���pM��K�8*C��K�1z�ӷ^�6�#��0B��1�%Aq�_jߚ�k���7U���cn�L�g�^J���R�X���]�7�)0���9TTI!$�ā�=� �����IO؃��c���fF�̜�;6�u����!_d9��w�C<b�W��`��|;==�����=���-w��K����҅KlZ�4�X�fK�;Ɇ/z}��B�y.��D�l�r�j�U�U�F5�G��������z]s�&������z�o��Kw՘1����?��l�ї��f/)���2��#�שd^��ȿ����A���!�Wlb��S��>�;4���X{=z�����f(��5HW'����\��� ���C�q�7�$���rK���@ݪB	g�4�cو�����]⸆�
��ƻ�p9yy�	։)����<�5JmI`gw��3���K��	�=�#U
�m�J�o�+��M߁�����^nNbU��U�1�d�z�I�&Ħ��/�$�����A��k�A�8�<Jd_�F��yBif"��*��?�Y��G
�;�]a1֧��3V��y{�y`�zj���diy�P�!��_O��V�K,(ceS����n`�.E�;��P�Nd������L�]	�:	��Jſw���/\a�b�ʅ�R�<�߱~�:˘�<�XTU��Q�
^\��z��}�j���F4r� ��J9����bq�� -wpp�(�U�l�捼�)�8��B�i�s��XB�5����,-�_�8܊�^َ7�Ґ|��a�9����D|�ڴ%e����Os-ˈ�k<���H"�s��)�^�M�vFKG�Ɛ����*����iP�gTmk�̆�j!�z$қ7ma�s���k|�\���#Q
�����b��.*0|�(�=��|�t�_�n�u_��X˃�Ւ��X�M3Ԙ�
$j0a����$�1�5ڐm����O��ɪ�\�K�j�m�JJ��UK{U4S��$D�=P9���Y�po�dg�{sK�A��&c��
��������y�d�Z���ӗi��Ħ�����u1j���
�4S�Z��)Ƈ�}�FӜ�~5N\���V��Isuˤ!�S��ߔG�`"����4u����0���;�׏�J$c�1��-��C���I�j�i�c����e��	���<E�1O:�*�$R6���?�� �_�����ʬ;�	���M�jw1g�:� ��h��Ď7�3�����2���0����EN����PS[K�s��jr�i>���*D*�惤�7�P��цX�}�2���8����~0p��g� ��������B�!���QV�����_|�+<'E^?�$��Ź��n�;��9I��K�r������|��la��ж�T�B��`��l���Hy�߇�/�Δ]���K��
/�޼Y�8KR�������׸u��k�'̵��M+�F�ᤏ_�Ӷ�������;�^kY����yf���J/�s���%Կ~+��@t~Y_{�OaQ������?��'���K�5�_@*f�8]OW��ؿ����mt��q�����ݎ��h��p����#���>�Im~@��.�
�Vf��:��C~�&��c#^4�B���Z��������qީp7����о�{��.@��F[K*�kC�v�w�c�S�U� ƅ+"=�����m@2�/&>l��NV3�m�c����y�.V�ɮ��Q��4�K�^"0����g��P���B���͌�`��0�P�� �x�w��$�OT�aut�
7�^�17 l۪1
g 9-Ē�-��]�5��9\C�X�S�m�*�*���t�_G���Pa�z��t=�&�z��z�p�W`��ޓ����c�O;ls�%\�6e��1k�h��-*K�H1m_�*K�9omp¤��O�o���s���:��@��Qm��[\��c䦫��r!2�sG�,j/�~é?�s�����u�LxV�Z;_�'�Wo�k��	�_{[��J:���q�ޓ>����� �a�hy�2u�[�:P�|���Jq��2��S>jy���r(�01�@Hv��uP�X�~M��%��]�ٚ��w�o��vXo>	l�Rm�k� "!#��o\}b^n�H<Yn����D���f��q3_iZ�V7Uy�������q�)��֔���d��N���4qnZ���9�����P"�A�@��KpQ���	���?гxb����ʟ6ߦ�|��L.����g��~��V���R��yOf�_�'Z�z���k
)�ܳl��s�8¢�w�V�{/Yq��
Ek�������g�؜~1�g΅P�>��&	�T�,P�;�8o@�L�%�j�bէ�}��ON����ܠ���il��8o�yHU	9�pf�f�`,UK�-JT���ji���� }i��s	�AH<o��������5ؚ�R+�X�����Hř�b��2!o��>1��n����cJ��8y����U�C&"	Z��Nѥ���#���P`�E�;߱�nq�V�U���3��V?�Q,�,�5�kj����g[�r.5PҔ�Xh���9;HPQ�^hՔ���F,��Xx1+<�!�T(�m�_4�&��b�� ����u���Z /�e*�SU���)L��Ǜ,C�TW�����:�gek?� 
{���v|o��l��-�^Fm\2�i�i5��.	չ:8(�u?���p3��+�\��sCd��dff-���<�~�k�ߔ�Ԭ���$.Ǉ�F�kz_$;�J�N��u ��Wh.��u�.,-T���'{�3���߸d(���,��> ��J�I(�2κy����X��&=��a�)��o�j�R�&C��朏�a�.;D5��
��#�ݖ|c{A�1.H� z}S냾NѼH	ݫb�}�}��>��R�>> �CW*�h����0V������P�y�|���XS�ݐ�K<���E�dB�YC���/��(������=�oBˢk(	���>պ�H#뿯g�t��#H]s� ���Xɜ��i��g$���Lc� �����(љrh+�'�b�-�F?�����o^J>�A�gq��h!,�]��Q��*�|�Z���K���->zτ����sqi�ii�^ȼ�����zBK�os���?c���ᬬRf]�57��.6��u��E�ء�n�]���Y�0��,�<o䮫���	��˘��C<F�,�,썊&_uxN
{c2uqIK[z'30�� >
����M&A�2@�<7*)B�s£\�#��@�{�Fd�u��8bF"�9��M�i�kQ}�ͬ��-�U,���>G�n�o�����N�6��C�1,�x&�8s���'K�&���y��1,g���uh�� ��'��������K��N�>�_��a��k3O����qW���Y��eO5�C�u�;�gNo���Z�ȱ(�_o2�w�Ѳd�3nX�o��1�5��-X���V)T��L�Y�_�LQvđM�Ǖ(�E�"�T�;�")�VX:�j٦��^�fZHQdD�=?��cH���V��Nl���,lt� P�Yt�]�!��Goo.�����䗕��`ֹ��'����W�C�k��)E�:'��F	{������1}���Z�&ӄ�O�z}���b�(L�]���+��l�Ͼ�;n�qeB�Bl�o�/_2lW���.�6Ht�����VphG��ȭϳ�2���� c�s����kB��ŠD�Q�p��˺�d�������q;���|����]|�=�9"��"2b���2�.�2����m�h�V�
�����aƂT��c	!���F�%H��� �j~n��&�����ғ�R#�h��G��^?7�ւr��?�`SpH��hP�uU�ee	ͪ!L�𫦦�K�#̝�`�L���zĀ���Ɛ`*T���6l��#Z������E��c8��0��yqtZ\^�f�ޒi��&�o�e�rPl��Ɵ��y������ o��/�-�B#�r��
&�j�:7n�Im�eg�G+��d�k�f�{	#i*��4W�1O	�ې."s�d����f��Y�	����~��}F�c�39��t�������l�B��^I=�LҊ3D9h��I	Z�oz��5f�[{zR9�l=0�>@/�uNs�Ķ�|S[\_�}X{ći�6�񕉑�0��3�/�I5U.AO$�S��2%������TQ_7k^��U�����1���T���$3$�ӥ���OZ=n���-u+a^t�l����mm����������o<\���֜�ݖ�s��+7烰����G@�s1��‶�TA��'=����fL+�%�L��Х�e���.�n��Py�Mq�r9MmM��3\털�N[;"�3e�#���T�!b��싹��t/~�Y�[[b�Q���Wn[$؉.�]W�+Yi�2^�T�[����ԎLp�3�8t�="�G���]}�卤)/J�i�Z��(oy�Pmb�;�#M��2�l�}�j���˨���lGݦ���^�I��O��J�cӽU�x�:	����n��ޠV�O]Nx8f^�pӇSeK'���X�O:=YR8ǁ	����݊H.��@��4lXc,*l���=?��<<4OT����	#e�2�^]�8ԿL��+�2ЭM��l�o��n�c�\��$��H"�:yzc$:�����QWb�կ�]$���v�֊
�$���~�߯�n�/
87#�N���EsB"��w�7�Ԓ�:�'R����n6؇�p ��������J����	ݵ�Pʉ��Fd�*��㼨#��_EH�0*`b%]F�$���G}L����Bg��P����I}_W^�N��@��"���~e���n
�ELQi��1���k��j^��}����06iˊ�͖5)�W�7��G�`ii������[�x.��/=�$+M�'�|VG���*z>��dt�ՁH�')[rA{�z�lq�A^�hZc��t�#~���4��[K�oLE,(M�}.·���4����:��!#�	!�_�m圾V��׈�����ӡ[6b�bv`a�r���t&j�Nɛ���`�[/��mL;a|F����j�&5dO��(]�R�$p�8`��O���	A��������l4r)��,��E�q�ֻ�bɣ�T�BM�W�@��.�^!>!^,�5������L�|�������R�hcLh�D܌:DЀͥ��J��QP|��\�o��4���.�z<x��ԗ��:;�G�#%��{����� �ެ�DŜ	���-�DAyfQ���&?���Գ�yg���Ck3���b���c,�;1N��'ü���f�w� ��q���\�]]��q�ʩB��y�5獫�3�߿X��Gu����_���p��k��/�:G�C�&������Kdg���N�X����]'n^8���G&�b���Z���V����(\B�|ŕ�Ё�D<Z�0d^Ga��������:����I%h�Slؐ�T,|���W�QQ�s��(ci����L)�Huw�^�Z��|?0������Ff��(C�@�F���ߢ���T�S�ݒfS⅏�dq��s��͛���Nɐ�^�H0�tܬ�g�<6��zmRǓ�Fvݏ�Cd��ߐs@	�J�?�򲂆�}�(姍\����Z���]]��E��(��U�2��ֿ.%�+q����."��yS&��tVWWK�Abs��Ҽ=^��(D=X�T����
S���R����^2��[+�9�a��nn�����e���z�Z.�_+��>]����N���(Y
�
E}�zQ�u�+ݯ�\aQ^2�lx��~�,�+���'*�*`�r���<bJ��m��Ѽ2Z�aB�U��%O
aѢ���numۚ�����Ӎ��`� 6�V��o����m��ii�Y���=EVKQI�B��E�3��"s2�R��/�����-!>� Mp೿�ԗנ����y����<�����4C����a�y�Ni/��M�.�z��۫�8��'��%�vJ�l7��=�;��"�呟wz��#��x>&7�[��]'
}>�6)�#X�$�@4|p�
�`1Ȝ���KVu�����}�3w���.�v�E���d�ܐ�����Z׹I����~��\Sp�&J� J����%�M���+��Ɠ޹�a���	��r��bi
b;�}X�TGY��ܙI��C�R����b�_�rPo�{UU��}��f]�w��&*j�!�%���գ���K���y�y�s�9���5!a�F� ����ngƤB+t͐r������R�ӳ��H��i�Ph�YVzX�����<��,����o<͍��5/�>�`䖹�`.M)�0��{��!S�K��O`R<���t��<�BY��=��Ta�O��.}��#g�qC�0ms\A*��Y��1���}t�^i17kڢy��`�H������^��#k�lQ歉I�����P'�	O���&-d�ڬu�HM:��W����`�N�ߗ�8l�L'���8C]���	��)Q;��TK�ңPGFF���f���B�6e��Åޢ�L ���y�2��ֆ��U��/:6�PhUK��r28���I����g���W{�Oޫi�5"*�#�c�2�����V-�y'#
�x�?���	h�7$ 7~^�)�m����~�>���E��ei��<���#v]`ȳ�RK���O�?���h�Ζ	�����d0n�������pE~�!"\��rmdl�]7{h-	�v�r�f���$>ux���颷ו�H������#�*���$'�Z�1_�<vaVU�o^,�}�[R��JQr�#�_�t$c��L�c05c�{���R��xֺ+7��,U���RS�:2�_���'�IΜE���:�c؄~�+����,qr>����
���у��T�[-c���&�n�P��Ļ��\�N!7�����;;��QZ�3�����mɦ�Dd��x;���?��bk
ǚw�c<-Ha���6�0-��ϟ��>����\�KQ)+�}�Tόv/�H����4j�q܌3��t���%��n.ٗ��З,�o���bt@��v|y���֞�@u{�FB�!ǻ7��U_ɑ|Y����,�[Sc�D��@���Q�OR��RL~�/�D���z��p�1�..5��A!-��V��Oe�gK-C��o
�����2p�"?�����Ʀ�����f#!(!��G.P�=S����.0�C�B�&�;l�hL�,&�hc?|��٩,+P6f��}��E+�-ji�|ɉ��`�g~7/|K����������{��Z9�T��ur��ec{%�*�u�@H��yv���7��9	����d\ۋ��0�W��M�4'R�q��H�2���#~�b����.؉�_��TȮ�W$Z;�W��6�^�F5�������L�G^�[�/Ȱ\�Q��G��Ť��O���Ҟ��
"�M�'������M���(��׮�I�ڌ'[(9�e�q�0����ol�;�T3-���7aܰn-3�4�n��X�P/���Z���o^톘#44C�p���N��,_|��Qz>�S�4���i�?�W�)%��8�yAʪ�?�ҧ�V�������8�m2�&JQ�e�	�����*��*X�ܮ�ϐ�M���y�ݩA�$�/�����g����S�
�CB=}��7�0����k��x��@����}�G�	@0ɺ�bU��epl�l*@���I\�d��OGb���Ʃ]�BC�ڭ`�N�;%�R���5���dmm�|�Jף&/'����ƒS�����ׯ_m�u[W��Ҵ���<���{���6j17���$�����v�����K�$A��;#RP��6�m��Epᷞ˓ՒP�צ�gP�,���,�8�><A��H&)7�������[FV��������3�ڕ��%gŧ������oQ�H�|��<�J9�����M	ZP��A��f�$r�˜����(1�W511��sC�'�����6{`xDH!�Dױ]l���F�*/a�e������wWo)�ia��dh�Cz�K����G���;���|�aRyl�)Z��dD�56��o�;������Q�v�}�K����ִ`��Qz�ȉ�2�I��^���^� �!����"V��_I� ��Z�����Sa�6�+���W��Boe���~�m"�݁ 2Y��W�GN(}O��t�����va/�\�x]�+��T䥌��y0����z�WC:ӬQ��K	{�)8}8l�h�`�l���R��졜(lTHJ��_i �q�	R ��������Y̰A�i�{��P��;[_YY�7�������Vx�v��@f�8)!�ǯ#`���虎�r"��4��N����p�&�)�J�-�-
�.�-9���;{|O1���/��lee�2���k�ݍ:&4%?�RQ�
ql��6\#0�aQh�'�<<<<�>��Q��ޣ�¡�Yv��Ȣ;��٘��P�����-�ͨȹ%�Ύq:����݂�=���1���m��A0��>o��Zz�XP���YҘ/��*��9��TN�1w.�c�d�E#��<��YN�a2:�F1>�Hw/�kJ�:#�:��~\�pĻ��^���c�06�q�H�#�?���ժhc����F�L8�k? Qk�̈���������P>k�K%������eJ,�0��5�&������7nl��{oQ�*�4i֟�$$z?�	E������h��d���"��F.�@1���ߝ4nw�Ĉ�ڱ�� %-}k��5�/{	n�wm\V����x-�Y���?NOMi���&%�����Xq/bP��x#��`�bN��\�p��h�6��"�^��p4��i EH�"�}؟-4t�m�Eפ!J��Ņ9 �!i�����i;�#M�>�[\0��8�^�x�G
�Y@�}�;�3ꆇ��X�ܽLp��N|T�u�g{��0k����a�]W�BVk��:ZtN�#�����:���*��A"�`???�}u�(sq�J&�Z9l��3_�����'5���Ӎ�_��$%C��)����2�uxq����%����2��Z�-*@ڽ���?U76BQZ�T�����6�1T��5�})�;8x`>���f���O��=6�Rz^��O�G�h�@�ґ!n��S�y�;��A.x�>E���Q�����8�9P?k�����Q���g�1-�a�i�&�)Y6����B4��%>�ǐ��s�*�J���j4xuQ��|vn^����'"Q�<���pF���w,��#��FN^~5��6��<����j���!��A���J����_²�❎����={L�-�Fm]���w�ЍVXC�z-��!�����dyyYZu�/�g(=q���D��=O�F��LK�n��;Ol8La���PZe��[p3�b4�OR6�֋����xZ�	a�v���d�՞��)d����3yR(���<�����t||��_V�GR�3�y�Y������P��**��3+�M���2��'~�寔�Փ����&:p��mq�X���.6W��5�R{8��1�t�,G<��D�Ē�����0O���?>����Tl޹��Ơ�F"Uܞ}L�徺���L��xXN��c�)*��gl��ba��36V�
�~}-�p�����ފZ#���
<��U�Ĳ��VWu���.2�G�|r��+���궼���ѱ#B�y�# O�JO�vƻ3w����*����8-��;�U�7a�rF;�<Z�+��F�\C���{���=�'%V��M+��.3J�1������������޿�������^��spp�����^y|��L`x[j�`�q��:�!a�l�[a�{�w�I�YwyU��aX�ݪ�|�����*��l�V���;���("�}m�.�^
�:�4�v��z�*���f����{e���o䭥`��k��Z�����d��#����g��������s@����x����i�Y&�07����`��h-z���X��c��#����R�1Q5����ۼ<Sx86=���n=啅KX&���6Ð=�}o<�{�"E�3,�4���*��*�+������[L�"��R�^ٖX��- �� *:6����#�����"~g��|JW�k�́��������J�@밐�)?�5�	4�,h	;���W�~��B�!|ck�0��p�D�o�R�'!2^�b���QL٬�_.��xЧ�MM��VZ@�o\���~��}�8���d���4i��Y��7�2�V)� �j#�K�u7LNC�5��ߐ��Hgljz��_CS�zm/_"<"�C3eR�)�G�����9`ؤ���b��?�FFF:664��[R�H�`��U�WA��_�1�j��;��ub�f�ؽ�S����A���T�f44�N4���q�2�_F�ʓ!N�������ٗE��E�^��������*���]}�� []�"�5`{���J��[O�ǧu���T%�mkr���yo�dŚ��w1���%��	����xtMqKI.��]��O����5qR��7[�v�/�j�^T��[t���S�z9}�P�����^~}:����)�pb��A�c{-S������VM�؆��<�Il��~�8�y9��6�=)�Ц݆�D))���Y�.{�4���Y�x�+�T7�oٮ�(���~�	�TR1$��a|������3�L8�ښ��G�Pe8){Tov+
�� #c�ܗA�B7j,mV�����멅-]o�p�����(ABDJ:RRZ�;�n?ߐ���u���]���W�R~	J�N���BEN�Xj�o��ʸ���J��}�d��qJ#���x�0j`{���L$�?������T����=���gX���&h9>������eo�?����\l�3ϭ�v ���V �ﷷ�<q�?%��^E��]�玜�H~ O���y��2�t��㣧B�Q\��b���w$��*02(/�uM]�i�7
�S��{�0��d(0�x�K��d&���z�ax�)��R:�%'�+��[\99�T~��������0	D7�=2�7b���'�M��me��|Ai�\��I6yv��oW�~�ƫV��^]y�Ⱥ2�Ay2��;�E���32Nmmm}�,�|�Kln���7k̪f5Utj�����R{���bן�;;;�ז���F\������{��z`��a��A� [�
�1��n�imJ���]�	�.t��v�:���Z,:BD��}��@(��@:���H
���d`�q�4..�~����uF*�=6�m�m�$B+�e�U�B[�^ݘ>���h��O�A�

C`�=�
���~�"�����Q�z������'�O���()��)8*��gg���տ�w�+��_@������!�8�ܩ���q��\�<�o�ΰV\������N*�55+�a�R�RY���ψ.MU|z�,m_/����p���I��T����|�px��!<cѣ��P��������N�UL���ΊF�u���=�cw�|B���_���?��=�VD�{�G9e�G?�'�E�D�������y�j�7GΞϱ�H��F��c_Xj�o���#c����.��X�(�f�R����`���YmBa௜�o[��������g=zb|���v�I�&�n�G
j��~��u���q��M4�[e׵�� Ml�p�
��E���&&.���l��i� ��a��}u��frr+�ʓ�#�o�|p������d=�Jn>\'�������r��pdG�OO`���\�CL�^_�<���/G~=*#�|���K1�������	CB���,����b����71y?��30�!o�-gZTXxH�d��S	tz�~�_���kh4(���w��6�ͮ��7dٖﰎn_h+�7����9Ӎv��-�i�:�*a 8�P�a�E�!�f������<�A�������`_�����<�i�MR4Ջ���i��ZZB�WB��$�;�x�����usE>�Edu֣ ���S [R��y����.�ޑk�D���lrP�0oڧ#1�l�=<ȶV VWK���z4�|~f��T%Az�}é@;4�i��k��b���*���{ޣ)��MD؄=9��Y>DF9֮n�0�|�'��8�M�'f��W`��}�0�JfU�aa�t9����ܚW���8�ԑ���$�G6��0𥁭��$�y^���67�@�;�x27d������Q*%0'Z�'.B? ��,8�����#�qn�����z�،���)Q�����1��`�[�"�����Ty% ����0S�������z����5�����'M�~D��?�����ð9c[ߘ9��\�-�^��&ҧ�F����<X拁Ȋ������[ZZ:�F� +�h�Ɲj����m�9-e�EY�S��=5�Lb���<����N���|���7N.��w��\Vv��"#�\��}�g�*�Upv���q�q\���~{�b�w�D�xÓ�ƃ4��c��[B����R�?�!�3l���"]z�ǿ����~"����PV���o�1�Im�w Jbl3��D��	����!V��(R����Hv�d���z����8�yтɡ�mHM��>LR_0k'hoonHQռ���o*urv���b���݁��glb��~���?&��ti�/ �pX%N�s�À���2�!�'u��H��)y[޸`a���l��|n�)�Wv�������:G''ρ��S(((�����GGG�u[L�g7@i]c��#{�4.?K����?`���X�������SE.`�[%b�[N��Y[;��^K[hM��"Bam:EF�e���A���������TW;�$0VOL(F.�X�4�3�s�%Ըx}}}X;o=+ �\��'v�%����}$ EÙ[ZVh��/��n6���U.@��Y��!�[� ��6<=���gDފ�"I;Ie��A��(2�HQIIKi~��`^�w�K�;c��nĺ�/�G���ቜh��J0 ����Ӓt ��B�OT�����G|7y
cj�Y>�������z-����2$��u�7�x��%'&_�����x��S8	A�ѐ ��f�m#]��g)���ˆ��>ã�w+�v��"�c��p�&Ѹp�I{U���ȩ���o�fo�5�Z�wS�>b yb��p�=�؎3���W�����L6hfxO���{��t� )n����*�I��fu�z��+�敏7G�Ξ��ÓKK��������S;ٌW�8�KT^����b����g=!�M��F*E��G��G��JJ��W��F��B~�/�ii=v`
���~^��$� ��Ňǉ��rfu<�3�^b�V>�	y�7_.�_�Օ�g|GDj��R�y	m���l�
IT_rN^�����á�!��a��xč�����o��*�A��!b�g�C2ay�w���x� ���E�P�,MN:�����H���..��74<���[�5�?���CS�C��x�%��}���n^����Ԏ/�`iZٔ�VSs>[�R)6�aNs�CT�#|m���7�
A�@�J����h¼8�����؟�y~�G�!-E�ښ�s�8;9EG�NN-66�(�j�
v�*p��S��nӪJ��L�ǹ�+�>	��,�J
B�hfP�V+�Qu0�y
q���m�|-t�����M1z��RC˯��)�6����"I``!"��,X��;����pV�/��;Yz=�%2{Uٺ��P+M/��ȟ	&��5.
���!��+!��z�W^��٠��CB�PSd�}�����6^n���xU�W��1e�Q�ƙs���ua
�`Y��7�Ԋt�Tܶ+w��5�/|p�dl��.��N������B5�ϠY� ~�M���(�z<�a�t��)��ϏqZ���	w�����HHu��I�J�q�`�+�q1�G^�1�D�]�[�bil*�>�d���!j�������p@�daf�	�:���aw�j���8г�޵�e�;=-�k"�x�l����w�F�˒��,�/�͛6"S8���������|�1�?�&,'GƇҹ�Y�-��,;��u���k>���җC�%ZRJ����#��� �foE�W��C�p�2�>.���,�����Vn�Fa�A���V�B :������޵{������(FY*���ѽ B�l^.��w s����2D���B��guXA�����KV׌���Ϣ���L^��	�,F�C`�`�puu�h�O��
!�/ \��I5hvII�&��ohs-4��噀+��'o0VI��U�v���oh}߱��3��E/Q��8���;�c�GG�D�XR�(���95G���c7�W��F.��ްP���$�E(�������i80y���Dck�c���-��+���&FP�ྒྷb�)A�����,�>%'�f�S�`��sڢ�o����̌.�C2��'~X�0�m~.M�9��(_��ϴ'�õ���G��l����ܦ*@����ӛ��g�:|�=�V�ux�J�T���F<2�;��厸����������9⣩�{\�жÇR����;d��.�j��g�׆~ݘ�6q�VZ\���k��,�G���e����:��|�=�y#�@^�ϟ/i�����`}��1z���$�ȑ����֌������D�nsMo�~�/�D�Cd�{�r��x��	��ӵ@�{ ���Z�{'?�ޞ|���͕ϲ3��\�&��J�Q���6z�ϷЊ!��8�ch_��I�~t]�81�<\`V�G̸/�h��O�v���4 a�n���8����RT
�8yU~�UZ�8>�#�/��R��p��j��y= �*F�"U8}��&���sC����V�7�>�����V���KD�!4l�벑-�I"z���Β.a|?�f�pp��>����T��u~q��Z[S�m�`z��O�7���y|~E�G����Iyppt�r�����Sr����tt+9��kSu��\����Je%GD3͵rB#y��w*v#>n�rz����R�!�\V��Ą�����p��o(خ+��v�W̜>E�5��￸������ٝ��yHeE)bbd�)*m�u�)U]�����FsbZ�~&q���������z��v��6<,�*�3j'�I8�5�孤8�`D�lM3;>�b#��9�i���R��5���|����r��18}4*�#V���*~� 22b�)�}�C��8~>����ܗ
r��߉	��c�U� �f�X���c:33�m�f6t��zv�8��Ԕ�������z�"�ju�~���NS�7m�(S������_m�-�uA�~�5[[;UUW�]�G6$�4
��=ģ�D�� JZ��u��m���R~.*���Q�KS�'p�gF`�`��Á���쬥K�v���+���;����u}%i�Aֽ&r��
[.�|%%�47t6ȓ�\k�����=�J���=�y�����<�/�����{�VYl{�_����R�ع`�ޛ�0��,��)�����*%e!@�V|�u�P�J��ü�Fs�g9���+;N^Ӡ�kƿ'ޯ|�{|a���h�����x4�a{�瑝��R2��Y����Q{���tj�!��H��a>Z55�[������B�<�m��Sɓ�F��L�Sr���kU�k�i�?�����^�܌t+�"���XB�
�ښ٘��&}��v�ƈ�,3$ L�4���/s
���}�f���d���7 � ���T�u��|OD�g+ !-'��I��4�Cf%�1� �:),���8�[��떊	�b�<e�����Dc��-!�
���A�禋-l��K��/��}�t�7�,+/���i�f��yriY�S���L�������pc֟����}|L�������v��f�J�"^��4�yC�R�ԥ9L�t��[�MMW��N1zP(�"�}DȾ�SPO\��upo���W��'*�k���"�NB�\�Pihh��Y��6��?�9�Ƞ#����暛������!Yi��7���q�cc;Bz��~Y-|F$�-V9��{���"?n]�z�����`6}��F���4���*��}~/
�5�1Jjg�M�_ug����q�"9"1H�"H�� ҍtww�H7H�H�]�904�]R���s��/��5/X�s���?�a�{�Ғ��Y�y��ll�&���-���d;��KJJ�'��-9KX��;B�t���/R�h�¨��D�o�89O�$��AC7�VV�gA"�0�%�h˕�1�ų��P��Uḿ��jl&hgk�z�--���4��grx2��9�y��-���!g��uv|����m8��*l�w���[�{#�9Q ��~ة N�L(��w��2,1�'����	д�[�ߨf��f�������)~*�<��A��:#��z�"���:5���*������@� �Y���6 �n%��ub%�ծ�	�A���ޑW+>r���9=�/���m���e�ÂP�㟦�����ч���z'D9@-����RN�@j�EEEo߾�a�Ҟ���JRw��@R8X�Pۦ旅��A��s1@�3�����'�����^kWF�o�U$4u=Ι!�����yv<����grDԛ[ej``�f<���f8��0ł�_/�d����DT`�C�Yb�s�/s�)H��FT9!�����X��A�ӎ`%.�� �5~���$���q�ؖ��� �[�o�[�7�QI/�;M�&���?WO��j��Jl444�i@6n }�����9����E�ÈGr��,Ps�� 7�����D�-f�V�L��k�yUL�탞��;��?<9���]����Q͆�g"��bɁ�<>�2<���$$�F�Dq0������3�=�E枼QȜ�VV>�vU=�:��!����b5W0kg��	�n���ݐ�0 L��z���
mϽ�F�:?�WopNG�r̾�����C�I�2����^M}oWN'�(mXp��4)����������b�G��w"Y��"��q��52\:�CSNe�U��|�� ��!'JI�pv�X�[J԰1.�A�'�w[[�Q,�=�����L��t=��6B��>��~W���~���w�E�KH�������R��_PC��b���JRR��	R%�T�%�������Q����X�$��a҈ z���� �JÙ��F����������~�����/|���j�E��s\j�*y��y�>��;,x�A�1��t�#���' u�/tr}��p�� �7�

C؀X�4�Q�6����˛Ų
�X`GE�ݩǬO߄��
��0�2���ˑ�tp��67�8<00PKp��������-��J�,����j�c�?@���JH�;"K:���Ͻ����ա�<����UuX���66�c�#}L��|n�0�@��p̫���I
�/�l^�pm��������.��r��o~�:r1OdRG�7&�����3YЧnzii�h�z�T�M���{||�C��gv-7�3�>��S__�Pi���ko|v�K�},���4e>�����	}vf�Ҥ���^U�%g��a��*؞@MYY����E�#*������Yd߯��\��x���Qa>BeGܫ��X��*��$T���O���;����đ�YD�n��Uޡ��
bR>�O-�n�J~�N�ۘ~�gEϐ�F�pBJ�'~�w'�~��漋u�a�B�l��g�`6ML78�0`�E�+-���n�|��3��*�ed0��^]S󜥼�$o0��V?G��p8��1��� ��B��z� �Tc�:ba��X����nE[�19��׍���޶�<:��$�ܓ
����JO�!(y�N�i�q��g�t��1hD؟[ t���0L�Ia�70�����3AA�+�G7��"��55�/z�* 0*���ǧ�ߴ����O������� ����MMWI���2�)t�y����^f
� ����_��^y�zR��}�a����qO���a"ME1��̴c
�!:��@���zAdZ!���ac��k���Ilz��7dV�4��	Y
�M�bw�� �6����1�"�~�h��4S2��cd�?�*؍��]NN�/�G�Տ��=��>,H�; HG���j���Rk��d�,@��lW2�H�[1��سui���C���ފ�ƚ�R�g�6))�#��KK���(zJ�f���S8,�����*����8�
L�_�p�=�M��N����{	�\�sT�w� EaV�g�n��t^z���kv�|B�myf�'���Y�(��ڇd�/;���=���C<~�������:M`ӫ�w㥞�sjՈ�M)Hw�r������7���{'<!��q���R���u;2�>���t@0{��d���2{{�A��t�#��x����l�˿9�H2�J铆UO-��0O=�u��0�Q^N�{�9}w�$�e�}�#��n�*����#�'�V�d�؀���Vp>���=�b-/eʻ6������շHr��N�ﳝ]C��ډ%ߓ!�L���8g[�gX&bȟ���Mn�>e}���c�5`�QR�
X8{�ˎe���v�Z���F�H�9=����ÞKcQv�
�l�7�^L@�^J�ͼ��nn��R,�������GK�=�eՙt�fg��mK���ˡ
���9ˈ�D-��ڼ�<�OK9O�!9+𕲲2��M�DJYaM힇����c\�ojh�5��\���� Zٱ��]L]���va0X�q^9�Q����~^,M)��	���R�;��
O�/(���jW�PX��q���^�"�: \��q��E\����j$�+:"��$�|_tM&���5�y|xM��[�|��
�*ӷ/Ǻ������Q���l�l>�?����50Th�z����(��/����^:B���5L�h��{�w���II;U���-��1oٌ�҃�N ����w��I��:�X���|��Q�`�"e���Լ�Ȇ(Ƭ �K|3�g�<C��~ݨ�\�睌�N���{��C�/2ѸX��t=����Kq�QA���r��c|���������>�8k
CϜ:�~�Z|-=W<�f�`��ʂ�۞������մ;
A�W��~,]{R���SF��~O�*S�h��H���A��&�[�C��"�0m���7��gvo����K�R�B=��sN��^�.��/ �C���&�7x7c����Yb@���"�g�Њq�ET�(�w��t�+��Z�cbb� ����SZ����,���AR������r�v*�A��=6e7�ˡ��1��7��Tlɕ ߄�;�s��f�����57k3��p:����^��
���텎��M�ߟ�A��ۭ�S쫚�t}�>�a��g�����;����������W���,)�'$��{�����#c�C6��3y!yl�ں~�]�R����
j��Fv��qΒ'-Q�w?o�H��J��������G�y�<�?���ǴJ͚Z�����n�&�=�_5�[&���m�T���9����A��-hF�'�j8�ӊ�𰬐Á����Ն��{�ڹ��������dh�&bKKK�I��矕Q�����} �S�yb� �aLí��iQV3X�qt�xAP{�01���%���dIYY�m�#
���?Q5�I�XCL�	Y
����z�~�m'�]��Kz{y0�ȯ �eB�h�B�L�쬣�#�ė����}�G0rMVV�J����-��Ͷ{7t\�]J>��b��P�����yw��o�{��2/lŀ�}X�����$�C6H�"��R���qcF�t����2��Y���9�ɳ��rI�޵���	�3����^Q\L�b�5#�qk�/��b4���ǧf���{�R�Q`��>���z�*E� �7�O~�*[E.Q�8ݴ��	@�-�ezvc�|8��n�1!x��C�Q
K����cz�h��\7d���L6��\E1�[����S2�?/�ƈM���BQ�<�I�������>`�^&���Ǻ�Z�����CĠn///K��s#���U�:���̴N��S��<�g����|U��yTY>L�e�Ԩ���Ia�S�/r�;�L'�����Ke��Q�lmn*2�k��S�����K�ܮ	�`���]d�]�_'�1<����W�r��>�,"l�S�m߈CU'a=LU����R�>�'�S��l�%�� ����"�@��sX� �v������λ���5eO\��I����t�t[����ˁ#K�?a���X����S8�����zfۣ��+66�g��$�+�8�J0�^��rM�I�!���!@H�2��7QP7E��� Ĉ���7�4����p=	��w�!ؑ��7�֞�+�W�Pqv�ϗ~�ο_3Q(���1~��amCqb��+��g���k��S�M�T��r(~��(��Mܹ��ov��Z{{�@D� ��'�%�ڿxܱ�V���{V��A�zݦ�5JEn񍅏թS�w�W	��K	=�pp��(h?�Zx6��Yk^}=�
�Fb�u�0
T'xtyi���b-z�ɛ���u&�����\�FR!�'`%[[ۦ)��F�۫�G]ϲ�Th'�Dy__����,T�j�����y?Q��ES�n��-���X�y���渴��ұ�z}gg���4D�-_��m��{��;)�0>�QΈ�ME�A��.��Yi�t��2����5??������Ȝ�UF~o��oQ���[1ÿ��b���E��x#�p��������^���nDn��ϡ�|���>~��KR戈��)k�ѧ+�j����x��N��nFvûk�+�	8��j����t�_�h�� ��A�`C?����:�C���߮li��+��|޹��ͼ�<��)�g�(�)Z���0-7��*XYX�;*�b�ME�͡��ԕ�}ƴ�]��Ȉ{�M��g9��1��	��fD�TMo )Yk������d���
�	����L���1�iԪ��Z���S����JG��ul5=?_ k8?m���3��:�ﱟ�vݲN�������il2��I {���� �^�4�A�n9����p�[�����2�2��?���Hn���QR��-��DǞ#ŕ9{ǔ��'��*�\+z�HOO�?L�74��߿����c>�,0u���s���	�`E�k�[i�kV9�!:ޓت�N(͐� ӫ�$���m���
������q����G��m�=��l���t��=����6$��oX+�������BU9��嬳�sş_����>7K �^0�K��-ڑ m�HL*A���\���{3�([���^�����ĳ 	{�%cV��-�?^��];H��Z����V0��mz�<��ɡh�J<�P�M�!wĺЦ�y1Y"���N���8���/xߊ���[����$� X&���F������4߉/���M[H�5�R~d&2u~>��H�6R��۴���O���G\��Y��)��lU��Q�"*����2��M%�>�n��ֈ���e�>M��sx��H��_k�Ǿ��3��E�+�("R�=�IY�I�s5������c��얖�gX����_\\�}2@h�~2�bI܍v�����w�"7�5���}�Fp��a㥇)�Z{d�c�P-�HY��5q��0�K��*��r(d�����SBb�q���G��0l�V��1��w�6ԍ'<^��Cg�&ҹη�YF���ҟ�9��l����^���7Ȓ 7RSS�G߽���_5G�)P��v�9����׬��}A���aE� �Vz~~��o�CmDi�<�oE�~�$E���
)Ĝ��
���X]fbf6��G��.K��XA��S���#ۿi�=������ˑ C�ת��^ئ�"���!���8��|�ݦ�q�Q��0&S���y4��X�#Yn��|��f6͠(U��Ԝx�h�^JT�[����uZ\������R��	2��:����_sA����6���j��yĒ�ū� �򞓀��]��1@�y#螝��
�K|ţ��DV����l$%��c��.��Leȟ0�5�����׳}��,�깥��`�|�I?�ETb����1��U�/Ԉ���E|�{�N|8��)�/���\+����@������r��d��D�Eu�2Q@j���?pP�ϡ�~	��]�yKXyEGՓ�.�99�V��_z���Ѵ}#�{Ƹ��F4RC]��g/#����sX��-+��?Ol��8�=���Ա�񣶎;� ?;^�I=L����>�L�JqX����ʐ�o�m�^ɯy����5���4�r�����bu�r��9����gĕ� ���x���1��T����k7�X<�ɌC��ߧF�U1�RA�p�{�b��zڗUAi��Ѹ���t�v����{��d���L�
�cg��t���g�Ȧ`,«���9�"���-[+���d����(SU@rC��a����H"M��������m�y�3����Џo��������z_����>v&"(��F�E�����{@a�+K�.0��䖤���Y2gf^���/:��v"|_}�zq�n9��
$���F��-�s�7���Y���iy�������ҭ����y��%[艊��y�r��_@|�s�z���<?�����|�=oVmM����(#�?��0>��d�e�</dm	�3��C�A{�ʵ�ck��q{�Ly����h�@!�d�A����LF>�$5>?^ԇr��rwG������e��q9vAN�X����j`�����u�fa�I�`�~�eC��j�����`���}���p����}���y��de@�63�Q5�55]M��D�' ��v��_,�ʊ���2�>*��nT̯�+�	���!�f�܄����m�e�f)�檥G�zB�$�Z̿t�Ϊ��8�Ͽ>-K�ILgr�^\G_#*�4	�%���2!-�����b���ӧ��Pyjcgݯ��h5T5�4�@�`1���o����|���:�Q�Ě娉�?����y̥���G�_̬��ڸ{t�a�d'�P�v~$O���cud��#O��&�������Y2��%�M�?��GR8��չt(.�	s���v��"����)��o�A3 �{�QCcj�WQ�sC��a:�^�~DG��E��*:�t���r��9J�U�@ۻ1
��g�di��I.�S���4�G�>�i�=?�d;�h����+\�������L��>��K�۽ea�"̼'�lX_�1y�.C�EP��F�ST{tO�	c5㘫��<�B��Rl_�݉����y��= �#3��*�7��B'�c��PZ��І+BEO�7t�.**�CD��!�3���7�ȃ*�}Ŏ"���"o��h��ϛ��?n2[A2��_H���&��jJ�A!��_�:|8"t�J��.��	�[�s��<���g�.X��Lx�컍���a�Kj{��90R���EM���#_�cN��Q�9@�Oc���sa��C[�V�p��<�r��=w���������~���ݬTT���
�4�1p_$&%��Y���A��ϔ���\2��H�ӟ�<�9TM���q런'�qQbM=��t1Xv/��x�n94	������ډE�z�\��7����KN��:ߖ��� 1B�)�I#�j��Ν��DDӷ}�⮢�ÎL`P��b����(��1�A����w��9���(��dh� �!s�Vu#3ga"t��>/�ʩ��U��vk�r�>�B���~[����i}�N���W$H2�jrR��S���~�O'����P��������Za���HSt7\���y���čM�LΔzؖ��.Op�H���%����S0%�y���l�w���#kN�:�j��il٨����Yj����	8� ��6ԍ�ϑ���D�_CW��r�L��ng��I4}�����Ou�?����k-"�d^�1��ˌ˃/��U�P"�
\�{0:6Q_�1�W<~���r������4�PHփ�huXy����rγ� r���T���6v�
 ����oA ��2�$��)��~�E���neA-Yp&T�(>����8}��b��B���zz2$�D5̾���KJ��(�@�����-&���cd)����&Ҹr�z+�U�V�po(�i�GfB㽤Mi�Ҫ�ŗ����mh7(���l,�yp�b����	y����'�ͽ�'�Q<��S�2-w8�Gd���m(�Z2�E���"@��-��v�!������LPQ�;1F���i�ױyk���g��ʩ�O؊��#���Ko.���9K�ʴ)����m���e�N#�\i����>M��~�I@D$?W��a���\=��������Ϣb�
~��5�z8S!*��yH���~yqG�?tn�d��A�eKl�A5Y8����fh�XSK8�D��=�C5Ͼx8��fx�*[E6��.O�eߦ���J(1+�]��&��i��F��;1��ׅ������� �&	6%?7އ�H���[�"GO�*'�έ��t����<�hv���ɩ���.g����v�Ã�L�_��i�yֳ��ݴ��`�kK����1�V��X��I���Zf�a�g7������e#A$����	�X�Tt��v��(|���+�7e ����2��t�:<���DF�����U�\�k�!I;��w�L�`���$p ��_śD{vl�Nj��؏��� e%��e[�{ �$[�1�WV�_T�V�(�K1��{�6x�:�6����#����d�nIʫ����e�k���ь��z'1�^�8h�x���	-��
*_���b��vZ���8+�����>P�Т�s��.���H�]<��� �������{n,����9�uM�l��KJQ��Bޣ`�j�^����F�Oq����2h
x�-�Aj^��)KcE�{�:o>���A?u

�h�/�*))�Y���I���J�(��8�%�0��>O�>;c�m��A�mU��b�َ��y�iN&�}�e,��[����!��(�����L�B����p(�����\oڢ�k�2LU���t�NǸ-�rF�<"�HC##Z�0v�_Pi�-�CnQ��r�А�y��BUEl���� �+����vy�fX 畹�1)����}z�*K�~5��r��������G�aX�=��Aˉ"�a�؞C�삦�&c��K]=���NbD��m¨BIX���𻚪�ġ����������:��L���S���G��|�I+��>^mU�	eU��{<����.e�0�&E�uNԎ��n7��i�.ōԯ�"��4��z���$����������hdR�Z�����}�w;S���A"qTМ->e-F`����Ox�!���jO`�M���5ߖ��r�Q���5��f˙r���%��?�����k�hAS��{F/?�������1��߿��խ��%k�;���F�W�J�Qת��j9��I+z�y*D\ ��-��>���wȽw�nPo�#��lI�~���7G��gZ�!L��hC0�څ�>gXn	"
: �ina��\�1��>��t��	�dQ�eS�s����J�2&&��˛�ʇ�V/�STV�"����?R�H�=<B��֬�1Q�xQd�>�_��8�����c�p��D"�}�¿�L�N�~�G|d"�7�_ ��{��謂��TL2�r.���=v!�U�a��NN���n����mZ�jZ�޶�#B�q+t��b�z�	�r����k>g�*#�>�Uʡ��wt���G:2����04Y׽b�P����6CLp��㭍v�Q�KK���Q���~�O�=K�J���o���N���^ߔ��iS�>�5y.9	��NݷO��ᚱ��4���������DoY>͌G����ѓ0D��쀲����Ok._��{�)*�-�����s�!KPU��#��dY�bl�*0���,�Pm�~򓬳ʗn�w���	`��C5ߣ�?�'ۙ:��Z
r=�EXt�c8B�c�.G�.Xb�0#|	��Y��H��r��d��壢A�澮�-C��x,��]�	%�tfE'�{��,����bml�����g��祗�z����Е����R>p	��Qr��155�/�����tH݃�3Rz78(66��&f�]����̦�E�pE���{�0d��8��2o�c�?��(Xƫn�=�D]��F��n�V^�|�
K.�	���ga'�/�r�[�V[�-"e����iôk�Qd�������>�ol̙����F� ��k����Btb6f}��u-�*9��&�:79�K��l�jC������0���&Omb~c�Z�Hwr/�T���5\z�� }z*�q��/��<e�(	��mfg����?����<��»)�-j𭸸8�$�V��{t��e��={
,?�{�U��bu`��ťMT�Qe���=:�s�z��R�=�퍰U���ARm�ye�Tu�6�q5��?CkY|�/#������Y(��x�:�R�����v���f�T�('7ɦ��oN�&�z�������'��& ¨�J�y���o����'꯯LD ��7��ji�2��%u=*>f�v���<R����;���ZW�ċ�t�����C��#H�Sz��湗#��x4�Td����ڀ*�y�F/V ��/�����^2��Ҥ(hY�?���Y��b�lC��:!���M։LV�m��" f��݀j��{ۻ�ʻ%�m �w���E�G�,
Y*%�Dt�ښ�W�Zw�)�S�q|��Z�},�ĵ��~S�_ǥ��3o��G�d]�\��U�|��us�ݖ�X��ô��K/D� �"��J{��I����`�RG�x�|X�nmm�,ƴ|�H����5lY�-�8a�c^s����.��S��^w�UĖ5)h��K�n������[)�;��v���sd[ �]( 2��ӷ§��S�(�x�W��@P�{z�W�$����T��p׸���2�'��_xxJ��vA�s��)*$B3����llĽb�	�h��̂mA� S�,^U�Ǝ7��������v�t,����(<��Ƃ���ʓ���ǽ���6�0����pzz�G�-�	�Y+3��#����4/�.Z�.�YBD��@��B�����L5z�
.	�H���xȤ�_�2z�sMVl��뒇�&1fȚ�!���6aG��*t��ҧ��f�.+WA�5�#�r�6����l2�q�����;>��Q]le�60�Y;��`b'eW1,�� ;ȏB��FP��=E�rY��Y�MB���o���aQ���}qY�S;ˉ��N`̓˃�O�g.xȋ�Eˋ^�����}��p�﯐��L><��Ԣ�Ã����|xFs�������5ȖT|6e�B�6+>�xo�q�E�:�"�V����peQ}R{��ɐ9Y��FbN/�V��nɓ}�P���w_��M�]Y�f��Z����g�[��H�H�Χ��42e��5-�G��T]Ϥ�������SQ9�<lR�BR��ZS���p��.�qYC9����nK��H�g p�H�������z����`��&YxP�b�5x��gV���u��^���G*%{�	�$4��*��ǩ����U+cHm�L����#~	��	C�E�ل4"H�d#���=��pw�/C��1O��5Ϝ�u}��n�{�])�*_[箫�>>W�� >�r�[z�����Q�g��Í�U܇3�b(7W vƭ^��3�ߣ9Y�ßɵ����=�xo�L�MָH�� G�����5�F��,�P�����S�Ҥo5�y���GJtt�6��s�~�3%%1��g��{�[��7]	�=��9�s�] ���O��� r�vh�}��I]��=v��$SJ˵��+8�����Qi�叹������)S潇)��Kn�O}��S�@��xvv�&j�ψ���|�lͥ;�;�<�F�u���LZ�0�L*��'��Ώ;Ŋ9��W�,�[���9���{QQ�Cl�}E�	W!fk/���z��j��hX%����LM����;�r�+W��ڠ7s��^_'ŭ���T�LD\���?�� �d�l5��C<|,����߬�Jm�GLdv|�d�kP|p��EEJE
?���{M�4)D����G�u_c}��#g����#c��k��ۇM���Ǥ�jDz&�Y�Bp�Ԓ��_��H!i<R+ �K�Sd]&�����zX9��<5"~�]4�r5�p��S�<"�N�2��s�t~ZS�.���<�2L������<Qx�H*����b�i@SU��`�P���>�k�l ���5���ⴌ�;upc���~�D�nh6\��kz��g���wD#=����t~^�&��Qj�_@�5�PF��#Gg]nlA��v�*��f�0H�g���ʹc�{i>����GSD�m�J*�*�r3j2J���;	%�ք� �O;񛁏m����c⢹`e�S	�&���ۻ��oK���t��nG3,.������Ĉ�X\��V�RҊ� ����{摤��
	��؈�eD�c��wS#�ieo33<<'���������=)���;L&��T���4�,}�4"f��R�b�!ĺ�-zEN�UA2Q<�� �nȥ��XzA��^n�q�Gc�H'�������� ,>�{~t_�4��ߧ8�#�Xs�;��h��r�����B�*��W�?�p�k&#[[�7'A��u��?S�T��n&�P�LX)t�1Bqx>�<�`q��$��p�}��VPЏ����;֑*n�f��/�%�����VH"U��+���/���h�r�����\6�m��iv.�'ls벞�>�$t�bGs�ċ���Ede�_lR{FQI��u�suյӝ�:c?�?<2B,G�#F�W}X���.��z;ի�>���&Q��ޣt�p1k��k>&�Ev�|�Aя��G�LQk�k��,�铊�u�$��@��>X-j�;�IY���Y��U�����B�tu���������/��?��U���Dvww>������y�3��<�"G�lm%���6��?: ����a�"Q�GA�*��Ѝ������:�P���(�qC���I��Z<=�-�ǉ} 3{��0�د�%��)��q�\���I�<�c�A{���%����>>���O�2�"��6�����l����8� �r����lH1%\)a!��e��л|�܁��Uu���aQ������H��%%���/9e�{S�VF4��r���ބ3��O%w���{��t�({zΒr�Ŀyܭ��m�*�'��7G��HM�O��z�m�X�B <�p��F*rs����\K\^�1�����k���OHL�?�L�y5�)4��c��C������ؤ7��z�/(��".������{9�+��6������c��50��"� 礒�/11��Pb���a`X��`@�.��b�~��D��q��PK   )_�XR�/�+ �/ /   images/74eaab8e-d748-4f44-9179-11cdc4bcdf9e.pngD{T��vpwwע�ݵE�n��=�w(^��;w)�w�/�{��d�gO��w�yfw�peEDBD  �"'+�
 @�  ��a�Wn1�����_�  ���7��ǿ���RZ�_�̜�Mnnn,���NƆ��,v�����  9@NRL�=�x�͝H}nc�d�𴽱�A�ɓAN6 ��b9����bla�j�~�8� /�M�=-[e�p��l��g��2�FS�Jg�"��c���A���y�cz���(<E0�8��0���>2r�/�yN��:�8���N�!i���<-:�s���\���)��1��w����?� �u���\$><D6f��F5t��;���9�(#�Vn$T�b~�U;�����x�J,���Bt���/(K�i�,�_�ޝE��*I}<��M�|�b��I�۰mʫ�}Vd������1�'�@9RT�}y�0�X@ci�M�(��(t����Nȹ�[$Ǆύ���?����;�2`��.���Q%K{0Ƅ ��Ö/�G�8*�ٜߎ���XT�w�IY�ȗ�"v����O��Nؾ2��a���:�I�G�k�Rx�1�@�	P��X�	�অ!��1X��9! 3��A��p;�$��8�� r�H��z3@���@��b��4'����W|c�\�S��rP���U`X먊|�.?��4��Q�ͳB��}@rO][D�WC�]���G������ݵ�2274����v��_[� �WAs��̔p`��ʭ���j#/��,7
%��A�h�OT�c
������R�6�*�*�u���K	�Q���;	 (U���b@�-���A��f����8�)R��$=��݁���Ħ�뻱�~�DD����:oڻv�&0ҳ��|�[��g�g�Ň �8A�j�!�V�Q�C-[�=ʫ�~��ѻ"����B/��f���u -�x������$Ն���H5ʺT�zl'�i�s�,�ob��X] 	A��g�ontZ"�I�.����vGt��ֲۦ��q����`^* C��(��Vu��(R2Ա��/T�(tb*��8a݈��]#}F�������@<��<y���x�iR؀�ڐZ~������B� Y5|�蒭��|�d_��(��FK˗�D������Ҧ[>�~���*��>5�>X��M���o������+NA�Md�d ��~נWs�i�2n��o/�o���w������9�C�'��������_>�"�f�|
��X��E�A)t�݃�]��г(�3v�6��^�$�G��~p����X�}��?�0���4��$��/��N���J��l�=�b��X�i!�4��`�L��210K��7��o��]�fmD��a<�}�/H�n���eK��awZl��3#��	��ذe��B�9��!��6��5p�p������DQ@�K����
�0a�⌮��N����t�K��Of�0�ߛ9��qv���C��܄OƔ=D0�d>E�)�˅�JƇ#��	��\U7'�H����^��Xsa���w��q��a��i>�6m�Y\u>�S��g)�,����ǯj ��$0h��E�([7�/g��;���V�"SV&(	�9X�EL?�4���ngk�RȽ���u
W�?��md��'m��J��T&���/��B�qg��S�{[��@Z�]y���>�8�Is��v$�j^���=%���-��~i��@�5��)˳c��(0Ko<��.�����~4����+˴�x茢��;��(nJ{�ͽ��Ňe�e%���n��=#xEë��I���]�d�\g�HKC���D���V�:�HX>��p1O��{TK ������(���Cd�F���s���A�+ �)���_��%��ܿ��W�
d�J~�ryz{{R�@o?�s�1�?���}XAc�z�����*	������Q&߻�����3���Xe�Z�'�A�omS�wԯ��ֈ��rF�)|������&y.��lLb�;�4=ue�!e��;z/��dJ�䧁�	,���=����7x7��l�ՓH�3_	p���<F?K �V�CM�������Iu�I��k��qzFg�}Mw���DD�94s�c�;�؏�a����c/4l�5�%�� ܨ���ǩ�z����G_�F�߶Hhuv����ѿM�{����U�dD���gᑕ����C.ޞ�ʲ�Raߥ� �l31b��a�ġ �u��D0�����N�|?cp�T�ź6�$A.���>�tr�r�=о�Wɷ)�0��Ƈl0�D�q������߁6u��y�T���p�w�>�ؙ��m�O����"I]�\#1���U�xI�x5� Y�p��~bw�$(���9�� 7x)�2�����v����������<m�MjG��Эz$-�G�,;d����x���B�p�{�:�)��'��}0���k�?8�8=#csK��+��6���0�㡇7�,�Tѿ�aR�Sa�\���-0���]|e�O���:'�G�-g����o����`�<Q; ."ze��Y��4	ywg%���H�x��gd�)��� d55يio���RW�%|���	$�u����G/vG���S�{|�;�K<����_�cX2��H�� $��+���n�b�'l&_��s�*�����g%��7�z�޿�0��n�K������왔n/|0ܾc]�f+[Q!"��wh�a$?,�_ɺ`5 %&j�<���|W�"�8eMol�Pn�f�4�z���2����knh�!�D��_�/{�>��~�J�� ��D�8������#��$mV�7����C?�a�����O�_�-��d�ɜ��!�fW�.`[�z�_�Ϲ��ޘ�3!��|��l��k�9��>}��z�O?��w�z���4~�Y<��3�������_滒��������p~+p��A&t�h��((��a�3��#�$O�a��H���|��J��Yt�U�sw��1>��j!ɼ��E^4=�%ҏ�Ѿ\�FQ�^7��XZdTi�&p�xOW~q��b�%��n�y���2+	,����a�+���F%;��q>��JicL� �vc��Śln��W2��\��S)f�]�˙���ՙ��2lLdl��~�l�?�(r�.r�g�Y����=���%3�Z僯�I��?Q����G~\�����	��Be<�.��h)��h���蓼���iˌw��;��F+DJ����/��ߩK� !XS���w���m�����/��؂�P��=s���V0�ȴɡ2��4؊�0I�3l���q�DI{G5��U�WY�'-VӐe�bwո=����z�T2��yu&&�ا��sNG����=��Ga��w�k���͑ 4��q�q/������7	v�S��"Z��D��0��XX>�Lg4�R��5�א��ӗj��-^:$�B�g3l����LD���irn� �o{�\�oS��5���v�!ck�6�>4�>�-i��7�<����0�(��/�3x��y����Q�d#."DKPPm$ýSNRKX�7ӏ˵����M�2�6���V��jаҷހ�	��imz�vZ��	�pɿSMԘ�Q1�SS���z�d>>�\.Y�"��T�s0���r�A��~q��{`u���K��:q{�����ߋ!l��&�a��&�8��&����L勵/1xIA�Ƌt/Z��:�	����08��c痌���F�g���vF~-�+�����m4ٌ!�6�G�;nmP�%��X���̶w8����}~A�jN��bw�(q�����i� ���#��Q�z����שּׂ����Ξ�'gg�iEN͜4�JS?���}Uy�I�C�C�7��yc�jb�B��x9���!7(L������Vg��g�Ńp܏ɾT�O;7&��%i1��|m^6�/�y�w���&w,3I�^�Ei��aJ��;�A�dW�K�>�!�[i;�ľx�XpN�ڃ����W8zCs���[��/�P
߻�EJ���6������ Z#-ϫG���>V���Q����
-�ʁ�������=��K�����_�bQ(!O�i�o�h��ivԇ=�(%���|��m-\����<� ��]z9����	�`�i�����o�=��=���ۼ��@ht�`t���8�t��˘���ԔQ�P�cA���VтS\K{�����HQ�������{����=O�����Ū���e�h����݀k�>a"fԙHaUG#��w^y��/jq�/22�DS��&�eP�sfR��0XF�jp��A.]f�=&�0Q��� �"I�Ϩ����a����6I���2��1pșg�#�>q��׷+z�Xl��E+�īӣ|f���\���[2����zX0����?��p5*J��c��%�#��A��]�pJ���B�BXJ��
�E�؟�B!A���?8�����Mg�ݳm�6�^*��'!��mL\�++�/OQ��G\��
т2;O��<w���tB,v&L'�O�"���4ONx�na�v[lq?�}�n{�֕����5��*����3�~�-$�{�5�I.�������W� Ҁ��r��ϿY�8�P��=��g!�j2�(�H�y�-,l��(CC�1�(��aA��� ��=i����q@˞�ai{���x���e[��¥Ow����7`S��:}��|6�fd���Ut��&���?�����eKK�1Bn�a��mWt��L3�'f����CjNYp6��u�Y��3��8����a��/���#0Dz��;�=w�HBJbsz(>����]��l�X��vB����HK��L-���)*�A{-t�x�3�������?��v�%��m�Y�u�^$���8	Ptn�?&�֥�:-ir��ԃ��j;F��U�^J�8!Bو�����u��Wo��\��� h����Zv�}ȁ�7�8N�����T�vT�.֐���K!�b�=x��:6����5ӗ��+��9�>���og��:���`�F��h��� ��X��
�l��b���,����_���䥃$�E�ۻ�n+܉����~|�����i'N�+QW�~|��ܴV[hp^4H{����q��6�ǔ�=$!~��Kw2��!��m{ԝ	�菡��}�e�b�����EM�������Obb{}B|,L��g��a�H���.4�e�}��`]憙E���u����7�
�;����IԪ���07�a9�ui�!�^�=��5�_۱m�����E�4}<�]���M�c/��u��3F�^&��~�"�w4��ƕ�u- ���%#��H_�
&bqH����	YK$=6�7-,6B�����1�5���k۸�^=������	s֍��I
�o��*�Rb�9�k�W%J�~�-�X����D�=m�1����2E�JV�,�����w��14���i0�W��W��=,:���5�h�}7N}�%�{=$ ]�ƏqS�������-l�GB�δ d+i�<�`��G�~�^*����uk��q֝��R.���9���X
v'�U�Qn9���+7�c��C�89�M�UDz��D�6R,X����v�b�H���K_���s;�^/Z�Srs����2�Km���0�k�q�TyX*U�	�5C�\d�|��3c�\b�4�C�]���$�gb�x�-q=R����'��uf:O����P�nP�H(]N<h�u�.�[sgyۜ��M���0Q�>J�Y��ǰ`dq�i�e����P��%#���-�ȏ�����Q\,�
��O�➴b<˹@�3��4"�}LgB�;xB�3
�2:?���
i�[��4�$21��M���W��G��-�f${��W�B[��1�7o7Ľ�'�uCd|��*ݎ;���Ҵ�\�C�gŻ؀^_Iy�"��@���{�;Z_9c���w_��� ��H�GG�V�Yh?=y��,��U5&9k�mőV����ގ��sa�`ӗ�z��~`��@�!c����d����Klq�E,�E�R3GX��X�+�N������Ӌ�mV�j����~;.,�/���N�8�_�'r��m�)`�&���X�G-a�E,��A��Ƒ�G2 o�Y��/�`ڝ�œ���)�؍y�"ox��n�9>��F�s�1a������0�|���S]<>��?��Z�'�l��1a�;���`��(ei�F�C>�ȚVMP`Կ����re?B+&;�m�vg�~<�-��W]$fzm ������x�"L�r���m,	�Hf�
��63�
� D���F/�� 2K50I�������Vn���Ph2j�V�F����������˜&Ҡ�$U���:}��X�ܑ��V��m̾����7G�D,$�+{Ӽ��:]ҳ������Wn%��ߪ۟r5��:c�|��n�顬S���٨�����0uv�����ƻ �㧕[k�O��T�u��W�l��w��͍oi����=2R	?��36ÿg���O�ߚ�B�t���z8���wΒJ].�^�:^���Y��B~f��/�,�SFX�������}�&"�&|�
��f��:Oi���Z��դ�yq�X�r%O������dЭ3����?&���UOj�~AE�͗��h�)?�:D�-�����#r衎c�'1�N��a"s^�g����2)�%
��Ʈ�9�(Z�L̹k�@R2l�[^?=�0��(�&i{ ����y)��wZ�4�#��k.DM�H�jP5���B쯎�͕�*���kD� �n5��u���"�b����a����=-?/�p���<2h���g��!���s��*�ENT�*wd����(	I c;A��/�B���;M�^R�t��ɺ���t������$V1Rϳ��FZ��Z�-���b)S�-tS�׶V����C'�w̝\H��Y�z����N�~�,gլ^��a�1�|HΎ��U��U�~9��h��!f����`d�n�=�C�J�^�5�G��DrF���2��j�hf�D�V.��1P��9�=v�Z�������K�?>��QK1��K���l�s5[غ�������IS[��-��
"{ӆ�y���	7WL��,T�c+���w#F�m8���0f�F�Ҭ���ǁ1��1��0i��R�oe���aFj������:.2���,�p�����^�gTO�Ql�͠�0pA�ڧޫn�N�|?(ڎ*G_t6�����8�R�"���;$�ٗI0���JȜ"��_<.�.��R�r�U�P,����	�?6����ǂ���r&4�Ե���R�N噇�֩.T/	�U���kl�~|�Q]�N�L����ו��G��y����{d�!���X.zd�
�P+�e�[�����g�!��L��_|MuX7L���Ǒ��O���2�^n�����w��Q�~�6��PF���������-�O�
r�t�xu\9rB}��^���U��ȱa�Y_
���>��si�=�"���D�c�h�Xt��T�ƅ���[�8	������Ҋ�
nۋ1�d�U�jS�Wsiڣ8�R���h�՗�|]JI�σ�����K�>�ƽ�壠�6z�T�ocG���o���>(T�o����
L�$T�1b���>�	���e�Rn�呾D�hh�2��E�)�r�Ö���
�����Ӯ�}�����������S+��
�=��e¸��n���J��H����&��ԅ�ڗ[�粡E}^]N���rP}�ܝwm;4���%�ٸ���k
�J${i@*�଱�o����Vd��aB���<t����!��Ƹ�j�R�]�\b��c��&xԯ�{_�º�w!pw[=`��;�\�Lj�}��7�d� D��`��Y�h������U5N�W�z���ב%�������e�ud�10� #b���	���6��	֏�j�����j�O��b�U���iF��@������@^8�P�}%�h�֫���5�h�6A'm/%y=�o6��B*&q���^�o^M��y��[�� �3�(��C�H�B�ܚ�[��/���)���XjHST������?�s"�xI�6��l��)��;�y���̬��!ve����(��O�C��ƻwăS��ΰ�&�~�3� u��o5<�������U��\������2$���?^f�.�@�j��nPP���&�^�;e|c���FT�C�Lc��?��,�q���}�~��-o���:րY���}w#G����F.�I�ܢ��X_�>�������;私�|�ⁱ�W����]޶n��Sh��؞�USR���R	�JF���kVvoB��ϑ������q~�m�/��bsoMM�n��m���0���9�O+h=�Dc(s���3"�y����R0#��j�?o�ʗ��q c.*����>��k>�B���;Jsj��K���hEޕ�>	�l���� t�n�7���"���ܢS
�z��>&��n�k��-�U��3�*���c}Kĭ�Y�#�����j�͗%z.Jv: ���8o�6������jڏ����T���>��d�l.Vwڅ�;Dc�w�__5��fe�X�0�ht����������1@�c�,�����8��F�]h�9�����[i_�.<ߘb3�g�TU���8��W�`�;,��
��r��Qp"�)������Q�ئ�fS�	�84�( ����Rd�М��`7��#;�U���kHS�O; c ^jah3��6����B �k�Y\R疗K����7����8�cH�e|>��׶�Ț[�z��Ǭ���R���m�.%�n�}m�vEs%�V�H�s[]-"��%�u���չMEs%�OD�e����eŨ�΄�Wc>�J��кdFfi�m%{Uh��$b��jjXh�������b.�,q���x�e��)4�'n�����^���I���8�zpI@)�Ͼd���ݔ�Դʘ����v��"�g������K����M=�
���2�j�7����Δ(3�_#����F�,�z,��n�qh{��y�GAm�;5�n�C ��!�Ēϟu�޼MY��x�����7�ٵ�eb�J�vr�Z
����@�\̋�6�Y8�i��4����N龀b���YIbo��>=���Ȳ��Qu����DrS��\������<�`��봡��d�o����<n	���.��̇��^��H�����#��/�W8b�W���m�jb����q�����I�Ax%��&��6Xsp+Kd6`�Q���y�GvF&����Q���3.�a��@2Q�T����bo4r/
�7����������z��@�"��2 M�9}�l!�鲥�������Ε���ʷm9�/]@�XϢ��-*#"ZI/�����
a��5Y����GB�3��ҚK��A~�}@\<���^�B�[K{�����R�����)!K�N[V-�0]02:fͬ���)���GQ�jG�e�T�/ӛ@�璫���/sK]�}�vn.H�����H5�].t;XX�mN&�Ѯ�cι2�Q>��N�'����y0$,�nR�C��M��]N�6	N�`�Her-�=d����vx���c���t�Ʀ@D^��=�a�cU���� ~nA��#�b)��']�Q���Q��K�8.���d����e�Ua����u�yt��k*DK�:�(S�(u��d_�n�y�Mx���L�n(3�a��W^/yr��� ��uG��<T%p-�/|'7�*3-�왓n��Vn���Ƌ�
�$)-�,L���F�^���n�K�?g��q��D��ϼ�<R������@��}3G�[��g�+��x[�"�Z�n�E�Q���EzD��EI��J�$��2xIGId]<]�`�e֕I�tq�hQ�W��( ��4`�tHF?�T"��p�?�@��Y
���3$H��7���U�_K��t02RB>-��iD��E�ڐ��r��Ҳ�C��������A��:M�$k��u�Ib8VWH��$�_*"����[���k�`�V�!K��H͐Ѯ�n���)T���w|�`�I�	$�i�(�H�vYC'ǥ6��\��Y꥙h#�R=$���� ��֚�0����,��Wl���Z��y?z���o+qp�� ͝v����7i��<�0lj���x�M[w���O�l��ץg�̂@�+��L��^�6.g�]xD:``�:�F��8�Z�'v�g�(H}^_�������@�����C	�ܞ�ћ����Ve'�}xeOZ��k-��(^�<~�<D�*_��c"I�%��pa�}�By�����q���N��Νc<����?ѐ)��D��������A���P��m���w��K��esy-���R>|p�V�@��n�)~@BT�L/;�R.�ښ�6X$f:}�  ��u�)`΂MH�-X�A%���Ue�W�G��8�_\��P�'��r���"V���X3"���Li�N�a�K.֗���H��47/�-7�C�w/_�<-j�8��U����1I[Oz s��(@=�]�Bh�%q����{�Y���a\_�  �OFt��c�2{"6(x�4��3����2�^��S�L]�!��v�B��I(�H��[~��(А�Q
�D��5�b����oM1�|��mmIgl��uK�ϩ4U�D�C�9NUd�t,CQM�ok\Hm�T�Q�A2#p��0��f(�Զ�vk�ٺN���O���p�q|����
t�/��2�p��n�tug[��W�n��o��2-�3��.r��2m���������l~Cpnh�Gl�*\�ˋ*s�,���#|r�<4�e�L��Ѫy�Lz\I����׋����_y0~~v�����I������z���a�C�U���d(�?��G�gA��ø��|��:5]U��s7�B��,��iz�bI&ͳ��v��/�&�É�,0oi\ެ^^~��f7'��[�:�lC�f��)��e��������-�.2Zʩe��v�p��<�K��D*�B�[z��BJv�:���P��j,���~�}�ߋ���gv����&!}�u�j-?<)����0�(1)Rԩ�9V����J���	�X���)V�,%�X��dm����a���`2����?�]����ˀ��]�'��ߐ{EY��(4�����V�/���#G�uk�e�z(y�v:p����y���(=��؁L��>�6>� g��Q7Op���U�������,
��ZG�\r�ȹɊ�3u5��'
p�'�h����S��Md O�M���#��:y�I�t5-~| �����,Y����s,}�M�4E��P<J^A�F��`G�SFU�̅ɬ�(I����N��v7��m�8U:���Ę\����2L_;J�����N�F��ķԹ 5�'��U�(>c*�ЋsR�%���~f��s�w�`l����:�P�_`���꟔�l��X���h�q���p�������*)��z�@�N�FQV����@�lcJFJΈ$i����@>~#��w&`�y���J$��D�;�(��!���W���D�J���4:-,�R���گȱ�~����c�On�����dC��"�^8R(Y����9Z�ҢG���+����A�˃z�q�\	W*zJW]eWߦC��+�iddB�S�:��ؾ{n^��Ѩ�WA(pyloNJ}۹�p��pǣ���3ȿ��%RM(�.�v [��N1����p��f ��7ğ��C4�����[K��0�T��uH���=���L��S®�t���p�g���/f�s�دH(!�bTC��V}�j�P��d�;���L���z��On�VY5O#&2�J���`��T��Fvi$n������|_�-�Ǐ[5�!�l�&����h���#�/寭U��l�DL��LXy�"�d��V�Q���S�=A`�cڴ��'՞ȅP��-�VL�N�����M��>m<I ���jFzn��'��[���RS|�b��2���ۚ䌲�f	8�mw~mф=����pi��R@��3�5Ԍ1���_L:�&^?�.�0�H`J�cL>I���G�֠��w[@_��'Zq.�W�/�c�bMg��繼 ���.����ra8��͹�C)Go��%�@l9��YgA�UI�]�?��\�It���͹�n����%ؘ0�+5,�Y�ڼ�g�	���q��[%��6���d��b�I���$�|z�D���]�4�A�A3�ٗ���ϺE�}�>��z��ؤ$`(?a�����p:L�>����)��i �4R��-����(�Jb���Z(4	���/��+��K�����=��Ŀ#���Q���C�޵BD�k�8_K7�Sp�bY*����]ؾ�E�F"����A.�_P(O���n�j�&�_�=� GҢz�co����F,����������̋;���m�Ђ��@��r���ky���n�{�>Y34&B�����SJNN��M�I�V�΋��*r{a�R_�?�����b����6T��ȱP���Dw���I~hJ{��XI'*LfXjmd�FB���\��rf��2ub=v/=z��O� � �R�fG�BB�h�v̟^c��N��< ��t��i.���Rٝ��O���'@��3��/��Y� O&�����ٔWz��[�l�
��|������w����	D9i�}�>:R����)�>(1�<�b��kR8�&Tc��@���t-�"l��-,���2��b��;���i c�m�".�5���h����$)Nl�Ʃ�<C�n*�	;���W�^�՚���֋�8�����N�#t�����u�
U5�7~:����k��#հ�������l�ޡ��u�)+ރJƌ>�t��^�>����L�22cj,1�"BR9y`e���SU��.�b�kWX���X4�Qc�2`IP`I���}�&��`&�#��&����T�k��bv6��}���ՑL�����1��AB���Y��ݜX�d>�Į��ǿ���H��#f�B�n`x%�xdZ�qOg�#
L�@����,p0��7}Tq��0�oϗ�<Fs�P��Z�2�a	����J�=g�y���bzo�,&�a�g�a�H��9�ӯm*�	� q��u��Z�Ǥ Hjѽ^tY-
��U)]d#&)��C�iA� FQȘm ���QC�EC���$�c���T�}���F'�L�%���	� kg������q��k���b�GQ"����?[�|���$,����<M����Y���du�nz�$�=wB�c@�1X�a_�	���7�ם�N����%;vMl�5^7��t����#ډ1���f}��XG�e;�\2HD�و<�«�z'tS6Ӽ��¶%3�O���n��+&��ds�:�g��H��f�P]���4��*������Krz�oϓx��ƞ�)�BO�3�����g����h�]�6? Љy��R<�(�'',����Z�{�^�ƿr7K�*�G&�@и�5���%6:��;E��� ���x�E�h.�m3>e<�=�P�x�II�N=݅"F��[`��LXe������vI<�8E(��l5tl��S%b����4,�=���>16��y�E��awc�'�jf���G#0����o�f�_�GU�F?�7_�x�dEi�V�mG0���'ki/&���*o�^�Vr�j�M�"UoA�鏫����p�yb�%JM
냄�rB�����$���ї�XdU����c#����ٹ�D1�{�S�KǒF��+�<��k��#�ƽ��W���!���Z&�j�A�e5�)���1Pُ�m/5�4������Јz�nPT�������Q���h�m�D����8����P��o�.~*׀;mz�+�w�[�2af�p�й�>��$h��X ���;^>epSo�a^
 `�m�����	�3�_jl9�M^n��C˺��E������e>�Gi�ʧ#�r���r��f���v|�>�#�d�p�Ɠ_岒������
��;��7�g4����HU����lC������7j�՝Lqo~#�x�Ryُ�����K�B�i�h����͋�Q<�u�+\4�`�;>�[�v�b%⋠��
�o��+l����z(M�k���X� .7e�k;i��!�� �,�}w���*�M�I/|Ƹ�U?���p-�X���ئ'D059";~8�	~�2�1��z	T�����AG����M`�ڈ�;��8˖ʯ�&Ͽnx~�����2f�.>�|8�n3�6���s(����{$q��u���o��;=1��w?��*�0�0h2�)�E^ �b���e�6-i�@U��m-��Gƨ�hW�{T\=W������5n;�=�`�n���W���`�{.�3?~�Od�� ��ȉ��Gšo�j�!=�g!_�Z�����vyЫP��|���A�PQ]7:�/�n)���Οu:�Ë%_�]QN��$E��`.�|P���e�������/F�+B�Ji�D��V�����Ĉ�y��i�_��l���]���O��Gz�V�����f�1R�H��a���Ȯ]s��ͻv��hqq<-.�w�#�o51��H�-�x�(�7'�U��H`m���s�s�dؑy���e	�?���f��cJ�Dz�]����c����S6�S��vș�8���S��<��J#�jl��}W}	[oS��j܎(Ñ����G�+�Ƀ��x�1c#��|j
�]�B�\�/��\��B��3yV��.��P�"���d�hbϢ雴Q��녈�O��Kv���äu  ��\�>a`��]�פ�2���~  ^\Ը����@q�f%�MwEfT�2I=	�X�XٜwP ظǒ}��2�	�#��jd��A�U�����\ǊvT'3o�44������| �B4�{���ut"oD*��c3|�%%���~@�F�c���Q��/�~z!�RX%���E-�<�g�p��v��.�������?n�O재ܵ�^ZC���Ќ�W��;gdf��_2a�	�p�\���I����Co�{�ڎ@�+�iU���=j����'��3���2������� um�C�ѣN��Fu���%��҂�K<������bԓ`d�Z�`
F�5��LX��q���qA��sW2���޵LOΌ!�w7!BO�ǎ^��I���]�$�^IR�S����������ؙ��M!�s�'É0#���g��ݒ��ɹ�����j��V4t)�G�� 6����A�9}nC��Li�3�A��7�Ńxj5��\f����,=I	F�U!��I�d��g74r�_�%��*�����B&W�$|j혒���70:�\�;���a��n6%o�|�^��`�e�5}U���W��ל�ߘPr�{�-�V�l�O Υ|`2�ا���f��)�n)C[��S ��1Z��K����(�v��h3�1������\��e�e�BS�J�/�����A�qYo��)��J��&�����s�־'ᆹ<�4��)��R79�"������	�Z_�d�%��g��bS��W��>���gm6�fqHA*�H(��
�űd(���@b��n/��U���$���l0�=�a"W�ν?x	�B�>���9j�D��Ick�[EI�$�9��ec���DL��9ߎ�?�]n�|2�-z��
��;-C��|����ߌג{����p��Gq�
�L����%!�=uQ"�k9p��˲r�i�N�r_tjd����٥Т򃘓�M����.��F5D�out�]t��8��<Ԙ�����z���{p��ah�@�LB����Kяk:����U��~ÁN9��J0l&���T{� <\Q�#�(���/1��#��+!�=�D��f�m���T��w��,0Zn�H/�R!�RqvQ�\������8�� ����Jy푽jb�� �O(�6&]!���7�X_�*���EN#rq �/B_��8����]�<�%d��j���$�����p��VM<
iX.���l_�����n+E�5Ș�}RH�۞�|i�����H��@f�ȇ�sm3P>+�"( �mU:bL��0p�gJ_�	Vq�}��#��t&�Lh��gy��	�]�ܼ?�K��u��by�&g���#����+�I!�]�LV�'>���Ti�E����=��o����#��d¤#<�)��>C#K�f��M����}���XKd�'Ao�I�۸��+Q���#�NQh�&k� �h���|e�#M�`Q�r]�����:�s��YKGT $�[=��|)}E8\�����@}0��E*�S	J�p#��>���w������� �=�O��ژ��ӗ�H��c�sI��f(W�6LAf�r��� �^���$�����dr�-�v�J��3�^L�(8tbՌ�k�S�Qc�&�cԍM~U�6�3[Ҋ�'�Kk��X.'��x��=v2ւk��,�H� Z���k��wf��谮q;:d�7�~�Y��Jֳ�ؚR���oN�Ϗn+���/��� ��l6Z�}�L\�6�_��
~�؈[ڔ-��3s���W��E*������l�r�+E��>L~���;e����+�↶vq���Nq/����Nqw��R\(��Z��Ŋ����>O��0$�K^�YQJ����
�Aq�4�We�p�%�0{�ω��	T]����vۅUh���z��(���f�k��pK%�ۏ�.�J f��Ĕߎ�ͿAP}�X���Y�w�#�^ы�E��J2[v֝6���mʝNKZ�*4T���_!D=1*}"�a��Ƹ�����N-t
Fv:�R<�?��ֱ��.4��,d����6���߽
G,X-�w6ݸ���+7UY���W�^6YSMy�u�n�Lq���I��EYGa�D@]��l�gfb$� Xu8�)d���l�vUkDGQJ�w��6��Eg�VRW�0����ϋy-]<G���GQ��姨�oZ����[���#���� ���M5��� �}x6����5� ù,���x�b���t���.C�R	G�P��S�q�%�_�^������p�un}�:�_�����6�@�� .�lڧ ����,�*���+Aݟ��ߠz+l��o���gk�#�L��}iO��c\\�Ԗ�F3(���0xY0�$Q0/u[�y&.��a <����C~&�zI-�����+���N���7��hÐRzMZ宋☛�;$�܉�?y����T�g����۾�N�k�Rvݮ݁�Bj�;ue�n�0�:��W�:�Ŗ}�״����l��"L����x�v��=\c�w���!����d�G��]�ڍ+�!%�gs���y����m��:k�1=g��Şj�$n?)!��3��:��A�7݆r��#J2T�9��A]J�2���X[t� �5�bQ���ua<�)�Kj���y��n���6��M��S]�#���r^�j�$yB>?���O�?���8������I�~Ҳ�IHf���e��0/�哢Ѯ{ff�P�ިMD���j5�!�"~��Fi�?���JOc�چn�Bɪ�B���i��kji��8Q��Ah�)�'���(@��������2c�׎�ݭ��G����ä$��>/�D�i��GEص�1w�����|��j���f������V���><QLB�1����\�Ѯ�c�G�dDJ����A���!r�:uPm{0��\����2����5��a��؃%'T��˹2B�B*mx�ޥc��.-��7���H����
s�˲#�Z�.��S".x#}	�i����Xp9�[�u��Pַ�Y��@t�4�P�!l*U3i�ɼ6��`_W��`ͻ��l���k٣�	󠥉[������>��w}���l5�e�pP`���"�q��B_w�uJ6)>t]������j�����nk���:c�``I�53���y2(X�mR�!kI;��ċ��l��q�)i�Qo�w�r����{��-	}�ʋY����v����Yvx^�����Ǖ�a�󕓟�ewGjk^W%��[
	 P��EH5��d�-�;W�G�9pд���#�<Z��m��R
/�g+���,��;C�	9��0�����5G <���4��S\�!���S.���Z�̂̓�ʠ��o=��ҡ���R�|؅aH�2�|�$��_k#�V{3�'s]�qǒ�x���c�1�?K���t�>�5��_�V)aϜ�=L�jq�����>��u/HBy��=���P�>�Dd;d5Gn�;z�.���isƜ9�J�=1f'��U�rB񄝆S*6��TdЫ~A췏ơ+{H�\������$ ym�X�Ȋ�7Sn���Z?]	v��V��hw�zE�\7U�a����Y7�������+�@��P�>"'4��؋%��� !p���>�H��,6s�`�q�C,0>�"��!/���l�4b xs�h�c=�썴^s���X�=%	���Ȣ?h���K����.��R�Y��n
�d�sK<DC��5���ھ���^��έ�D���_�Q�ίx+�=ՐN����Y�G�Y>���uZ�W��Y�}�mݾ��?�w��p��,�Z�^����ܶ[S_�[<�w�N�ff�����B1d����:���C���2��{��䦇o��'����Z�r�Zǜ�&&�ɮO�V�l������p����RJ��oU(�JŎ��yfY�X�gm;�"~�7��N*����,�T!��X��;��F�+v/������9��#?q[?/��{lD����o��?�౴���W�ִ[�|���d�)�~�{w����w!sFw�̆3�4����ԲR�`���*
;�,���X��ܵ"��m&d�:t�2c(T�	:� _�Ag�_K���W�D�'�'�.�D����E�l�G�^��x��~�vq��Rc��ohF_U����0<B��Xb.���0��
��X)2�˪�a" ]K>q�,��9�	F9�og!	z��	
P���]s�i�A��|N�1%��46�RL����#g9��%:��[!z'��coNS,+9Q �L����òi���(l#{1~-.(�P��y>>B�}"�#P���6���Ӌ�7<�덷Dll��NAA��P]�I�,�NY��}�.wc2\��E�!�>|k��v	g��_���"����kuK��X��C�G�<���M�q��l�Tz0�1`���L��<��B���/z�~�h�~2:~-��X ��:�a;v����j���wL(���%�23��ϲ��yZ��cT�Q��:/||/Racݧ��їb3�.?�A7�I��)��@[r�,
n�	�=�"?VpR/<�n@䉩��D�����7=f|��1�Q�_rmA��x�T}��F����ӂ/J BJjc�����\�;��n�
ȹ���������d�R��U���,����67-�)m�DW�7K�tM�Q��;u(a�eb7׎�y�I;O[6f�U���	�;d&B(Q)c�i|<d�����6�����IWgqY2����І��˕���:#'I�h\��I��:��xI��3\��-��_����imo�(b�hE�`Oy�㡃jц�����K���N��v�R��2E��ޓ��|Lp_�n�c]��7�bp��Q���5��G=���]�>���q�,����+{�W�O��Y(+W�Ge�Y���c���+Ne�'
~�Z���ru~��wK�[t��!�3CR:6$122.�(�!��"h�.R[ƏU��[+���{��),n=߹�]�Ʌ�L����ʩ�6dɯr�b��m_�TΖ6*C#+8�k�ި�Će�� ݸc�PzU�����X�p�"�&{�T����bkԹ��� T49�}��ا���?��}�+�K$\�"�Itg,�#�L�/N��v���0�fc)�h)������I���������}{ޗN��,3sb�ݪ�񰝞��+d/�vZ(ެ�+dC�����cU�ܙ3��j6�n��)�VV:��R�]� ��~(dZ���f�.����۪O�����w�c�7��!HPd�&�v:��P��m�f��R�^��]�Cf|6ܿ�F�#ސ"����lTFa����%���9[�~Ҵ,Xon6���,:D��e�K{�#�j�09�R뜓�D���t+�{���?�дZ�U�����<���CW𾷒�\��ٷ��]Tn63t�7��܋�LʓF��!5"�DB�-5�֐�a�0�f$M�_�*)��Vs�=�<9C���m+�1�[�������w�h�=C�C�f�
4����N��#�	��b"w~ht��x��Hi�6V�r�|�4�O$3M6���c�p|� ��@ �z�f�z6u0D�V�FĜ��渳����|m�X/�ӐKG��"���4�8��W��Gi���FO�]0o%��}N����ֶ	�Dt���Y�EW�ڙ����:�������Şw��}��~�A�K�������qK�)g���j�L%|��.���Q��v�;�T�G2B�Yh����:ߠ/�����p)�%��U�U�ɢ��$.�L4�w �~[ǆ���>x��״H�`n�3�{x��>9`6{�ӟj#;�+;�d�"����FH��9�ۺE�Q[#�m�WŬѷUr��ǍUZ�Ә�	�5� =/�~���tY�q����~� ��+D�*59������|C	[���PN�P�{o���⮘��g+I�_H������m��=b�%&��p<V�	$��;q�g�جH�O��6�el�L%U��iF�v[�6��޻qh	P�FɅ�z���H��I�|_WvRc!h�=��U��Q���}	�~6���D�kC�Or�b���Z��i�~��V��+��wTn���e����]>��G����\|8XM��ϻ�d��D BG
9��������,��:^CR�<H����Ӯ#3V��$O��tւ�j��U�Qa����ݏ����U� �V�xF5�J�c��
5��n��4m��cXR�|Q�0�7���R�[7rkͱ8O|���ߔ�0ζ��X?-4X���1�M�"�֗ �t��`/Wwt&F��[�v)���	�>�Uv�͈���Ѵm�������o0O<����r������ڈ<�e���Y�K��K7C��Ұ�r��oM�TAW�]<S� �iZB<����l�{^��p�XtR�Y�?��ʡ��牢����8Єǫ6A���Hs�����ѝ|�D@��R��T¡���od�� ^�_��x��*!Ǭ��+�v�������LK����uer%�Hz��?u��NX�[f9�_\9��m�䙪ֳo�s�NnT{��K���l)�uSZJ�(���׻�	��c/>XEO��4�dS&'
��}6��kF�����OT���5��f��S�FahH��p��YO��g���>v*6�C�[�@��l��'�pQ���B��C��M���1�����2'�خ��t�'���®�q( �Q�HRǏ�(�Ӌ��I �o��pr$��i��$�[��e����!����8��
��[��f|�)�)@(m6���2���S=��q4�f�G]}��	���q�^k�����e�H?ub2;yH~�g!���(��'<Ia�>��X�)un�S���Ac�O��4R,�H��~����/f.Wbs4��{���P��/�����O� a��q�=� ����Z�s�ĲUu�WDJ��ݶ��0#���_J�s��)�'���ZCY(H�>���ߚe�GE�Ђ*a�$j
��8��E(غ���S��n�x��i�z�ꀐ��1�A}^
�Ѭ?�ۯ����^S��xS�<A4����"��B���ѻ���e�3Oǌ��t5��Hڥ;�Sf�U͈�<VK��3#Ӌ���z-r>ו*�^d���5��Z�n�.��[�ő���Q^m��ǀ�E�P��M�&F��CQ	!���,�	V��7
t��sh�JLY�-$��Yx����|�z��K��,̱�>|�2�n�˒�[�y|��n+�å�=�6{�F,��t��G�8���8�Z\2�V�Vƈ��O�5508�T��D�ȋ�3I��H-E�-c
�x8/�	բ4��H��[	��!�'��դ��� {�ehD���8��;"<&����R�y����P�D�1"G����q��Y.׊�7F?�fb���{R9\��}�x�����v
4�-���Q=E$D�e1j �e|�;9���%8j�x���,�9
�;ev�� �mԳ
�a�3�O����Y�1ZLQ�
�hL;z埄]3v4�Dz��"
 � 3bW��DO���lZ��ת#�`�c��y�R��Q��+���M���dC����u�m)����ұf�m4��ݗ:���	]H��:a�ȩ+W�L[����a���49N�~s_�v�c���Z��[�u��/>�y^�Rf�g��V7S��H�e/�T~r����E/��s�o�i:Wƾ�SHZo��Խr��J�ae2�w��s���SP�ß{ԩ����v�O#=�]V�}��(71�O�kb�m:�=c�ۼ�H�ǶغEsﰘֶO��,v�֍7�-�3"B�ɨ~B^^�"Խ�x$�+�b���i�q#S+��P ����� d�˰��;?�ڥ��Zrj�?N�.�q~b�!Mp��\�V����+j��;�9�5�\-0l�c��!]ɩh�&$�g��Ԥ�7Mrl;��.}��3%��=��
 &��-|1�vG����
�K��2�����V�X+ᧄ,?���Lc��U�Z�6w?�.�p��w[�i	��Fc�sfV�j��9��C^��π�j�l"Y������B��.���#-��4V������u��`F�b�*��*�6��a�8د��Z���I������a����u�*R�ƍ�R�(/�i���5z��?`�v���"�2U�����IU��յғ"�cgjЀa���C5{�s��R^vf��Yc�\��.�����(�[H�� �ӵ���F��o�w��@2w��J�1��̤���2Ӕ��H�e{sv�<��Er��>���e@�3%���ǑPˡj�p2���
9�͚�WiA��>Ĵ�4�#��喂1t�Ԟ�<�C���>ҝ��P��U���O�I�c����H�KBa�vOp���T �>8W�c� d�gw>���!C��K�Av�²!���Ȃ�Y����������;I��&���Z��y{o�l�Ջ��<�+�ܷK����	��	Nv��h�Q�@)D�,شWW�v����CQ{�>S>��[l�Bi��p!;�}Et��1���Ką����Q�����3����ks-в`�d�Ȧ�Z>�F����fws�M��.����w�9/._���o�Z�78x1ZX�8]��Bj�\�5vu�'�_�7���ŶyhE��k�����ϸ�e�9`O�ڝ����o	�>��j��DF�3�}�b����WKf�m-��}���͵Z��� .vZz՝'��D�q���O�|�3�x����`�R��?1�T�1�X@o�c�W���ƴ������0s�i�C8��;�� ���#��J����v;�·��E6:,�\G��6x��Ȯ4��E�����D}*���9@���ǓF�e����Y����g#P^�͞�W{8H�^���b|�,�aL9	��UA���ZG�pH��#�y�w7�bU�D}��LFX�T�gk`��L�K	"n��M������p�cc%*�Jn2⒬ʇ15��+W��� �>-P��V}ܛ�� ��i}?ME�����ӛ�vd(1��&� �Zn�N�MW�賕4m�.0�(�E���<j)��b.�&�aTf+��`�t��맋@���d��5��3#.���q�� ��g�Wy<�X���Ch?�`��xc�QJUMǒ��}z�H}��b����M�gm�rB��?��|$a02_~(�ɟ][d��m��.U��KOI>���]�����ҥXJ�������P��0<�bՄ��f�A\�Zg{�f�Q0��:׾�{���C�;���G�媹R�q�s�n������B[��54v�)�뼝*�:��^�~�ZQ��5�$�&���W<R}��U�dC�?��V��oM{-=��9�����¬�Z���| ����`'?�d�*�:d~�xl,Dިi�Pn7���9�Gm8�S;��C$+sҀ�B��`�@d}�%d��zIYyĂ¸?1V��Q�Z%jpPOP��~��i��7�vO�(����k�	.�(;�uIÿ��ʥ�b���ge�b���pD^AK�'�kI"n����'a�B��"=��c��Ȯ=.�h7F5s��P�r[Γ2�A��y���QnaPJ���?��W��}Ҟ�m�%�Qjiq��df��{U��DH��W6��y����5Ŗ�~��������CKܒ�[�k�w
�z���L�\�Fii�k������_�qW�����W��`��� ��eC���5�mY]�����M������� �&J�>5g-�|�(E
9�`+?Q�tu�
���G��1�=���3�1x���rޯ��~�0���%����\�}�y{�'�i ���fgV�!p�ߋ�+J(�;��3��~��/}@��l��L^rD58����zc��}�v��X�\�*�r����T���iy?�	�$V�9z���ػ�jdD[�YY����`�D����vL�F�
z�ǁ�f�:��R�F���!�np$PO{���+��@'����q��M���:���������ʖ��Yi����B�q������Y�K&�LEZ⤃�L���*�%�����QzY� E������?��6����q�%�ɏB*�-�s�թ��KQ�v*[=��O�/Zb��f�/��J�[(��C3��?<'���� ,6:i� �jً���F��i{©���Fs��W!��/l�F�j8H ²�q1&�y�"�k��f ��H�	�Y��TuD�I�5~�z�ĝE*f�P@a�����V�٧�� �\���"b�%\�!�����R���[+�ˆ��ڹ �Bn��cw��I�7����{��t�A`�=r�-R�R���3��XؘV�B��Lz�T���u�������\�SUȜQѸ0Ч�ϫm|8 z=[ی�Ը�]�"ty���4OH����g_\�6v#\��`Ț�c%ow�I���A����zj��������L�Y����g3>�5Y��!�|5"��R���[U+������ŀ��Qr�~U�Z&�3��a�Ak�:#��I�k�*����n���)� U�J�g�>�����^���q3�A�HH�{i�ެ
9�!;�n��S�Jͥ�d�Ř�,�C�k�k�KV;Q��pB�(1L`�� �9�+��|�ː�q�Y���އ�k�� s����=�Q��-�`��T(I[��F	چ(�޹�׾���7�)h9d���E�&����0�L�C�|�������|��@�㄂wrXҨ�;wi�����b�b����28�`�R�&8��-�,����6B��+EZ��a�O�|G.g��dm�j��srFn�1����HP*��aM���O�R��`6�Jk���K� �l�AW�;"b2J���<pT�%�X��Ua�A4@�|Ɯ�G��;�k�g��t�+g>���?;�����Zr\	����Q��n�o�F& @�<��P瓬�wUw	p��u�-7�¬�x�ق֢��p����!�*�����n5�J��@�5A��%p�gW��u���W1���X�/G���#&����.@9�F��!�����ռ�`�� �Z�]커o݄;�ȑ`���c 7v������6Ԣc9f�b�����Rw������i��mJ/.�/���4?F�0�z��D����olO瞌,T�1-K`��R�H%tb��@����2>��8�tmB������Mj�C$��Țn�O���k��Fz4���2��c��{6wX6}��n���X)co�����Gr"�� g�S$���Đ��1�S�<���0z��v����K��o���~��_��v�b�$x�XY�1�����Y�]=hk&�8��99@�w	�Ovz~"��Ak�xoƢr��ҙtG��2|�8�4�[n��7X�rЭ�T����~�CM��� �}n_�Ό����W�� �%|���/ӻ�L��L!d=�u�+D|���xQ�����JN$$����I-�`���]_�
��c[hڐ�w|��q�$�����[�E
�:���}?0[�.��c�Ѩ��"���ɖ�T	=R=���6�����Z�'�?i������]���2�;F#������\�����.|�F��:.9�D��!·<�n*	tY��0���l:]Mݢ�#�0�x~���^���r��o�c"g	�c&z
.W�G7��M\�^���o��}�r�������}�blHߟ� ��y�4n����4�0�raL��Ur������#�Q�^�b�\���
{�P�]����I�U��R����9�.�>)A�Eם����9�ѱ4%m���,F=k���ŀ��|
"�0wߕ�]����o4��wn:�J#�XL��>$�%$�8�I��'?�L�'��J�k��5�!�^�}v�MG2ZX�9}�i��_�G9��Z��ԭ�'�uχm�O��Z;��s����+�m�2�祚���7���k�ZF�����C�t����R��C���!�]��^�.7`5ol�h�C;�0�_���3�(��&Q���βR-�	'(��3����T��"i���GS������V~�g�8u�u���N}c�	�=N�_RJs}"[y{j�P�r��C�����oG�E�{��N�����$b�CLм�B1d������ii���ќ������J�e6N�0�!y&F��Ew�H!�ب�K^�4Q�6�&��H-�6z(�[���4N���밅le��^O��T�(E|4I�&1D��ShЗ��g�I���W�P��F������2�qw�\��Z���}ޅ6:��%A���EܥA¦a������.ʈq�GX��˞��Im�1/ץ��/r��j�m��i?�m0��$!�t��ʁ�w]X/|'��ע_���[-V��w6��/����o��br�,�J$t���s&�o(�J��
���>�����RA@�Ƈ�^���ܧ��d�t�9��?S`��������y6��WZ1�l	}d4��-�!ˏ�2z����z�3)E�<X��}�;Fb7V @RW�{�h��_��bӿ?,����G$����;�w�wV�T�li���e�_�� �����`��3c��[q b��~R����+&l#-��4����+>���l[��B��콦�WFU��8�=;�~΅��O	��6MZQ*�\�G|n�E��������.���'�����^��Eܡ���3�vF��7����{Ý["_����(���u�Ŝr�>�Xk2�ܔ2��dq񶻇Y(J%����j|۶��t��m��d�v�C+�^ٗm�'�?� ��6�a5��˶��>y3�Ie����v+5�Y�?��o�}�� ��Eޮ�1�Ƿ\���O��o�����D���,a�����Ih۩�B��#ţ�_T�AӺ�L�cU����/�\g }��� +c���@(m֐žė7n)A�>����A�od�����B+=��烪U�nC��
�(zZ�$v���L�ˮ��yxG!��Ga���kw�T�u�!
OZLLI{{���P�PB��_q��}�EA�s��d��ʙ�żЕ�5ѥ�sO2{�J��m$P?ބ�$}��	��y+�yu���5�jF����
��X�&H���é�����-��` w�]���&[�}�h ���<T΄��qԊ��9<Ū��lm��@L�A
�8υ�~`Ef��ZsV�_�~��|ԗ.UR4�U��Ƅ=�"B��J��"V~� �+굸"�D��q����L����R��Zh��7�}��I�r�r�l>�U@u�l��@��J�b��yy)և����h�ՆQ��#�Ұ"��7�֝a�rd.���Q�{?/ٓvc��* ��<�Jt�RW��f��]���|'<��/Nx����L���_��0�<��¯��K�\�E�c)O��$G"�`�{K�ZR�<��ۣ�y��d��Y]E�CyH�ڒx��
)5�0�����nU�dy�m�H>�Z�S��N����l�UQ)cA�LhCh�G�>>�}>4CkZ�7�A�(R�,Z�8T� $�IȬ���$=.�#-<1����C������_��&�mk=
������}��vG���ˏ����JĪaeX`o9����j�v|l�V�h��vx���� 1~3\�.�Q{W�b�KMŪ�n�����ʂu;	��?�0b�$�STU-�|,A��r��
4�%e�)��b�P���BPiS!�9�V�w}{4��)�o�Q���1-��?E�m�����2�\�Gg��P��}
���V,f�<fa�=�-�RuG��{�쁂?-`)��Be]^�-:C�a�랕��IU��l�Ea��ʗ��F���Z~�>����B��Y�.Ϳ����r%��L^^) wC����m����Q��#�1v�uC���-�H53���-������N�-��ޙ,y��J&�56��H$WO߆	.fQ�.��LWm,��ݗ�����B�:=���Ь�mx�[��vo@�p����j|k�^��.�VveN���T�sayN�/�ԅ���H!>��]ip�Z ��ʯ0bx��5ZC���.F��{.U'?���Ie�T�\�,��/���s�tځ�оެ�%i՝C6�`pR�&Q�ېryq����M�Ä��,y�Cf�gߖ�+p.v�� g��8_p��0�mr�ic;��
|�^�ƹTȻ�Ub�뫝��up1'DI����˜D�s����^���"�/�&���tW+{��9�%�"�����e���=�a��1J蕕2��{�K`"�?�=1u�Bk9Q������u�S�$���8=���uvE	�E99����w��:3����g'�$����g��S�G����v�Jz���C�k�uo����%����J�J�}_b$d�t0y)oX��ȅ~F�wP���3I��l�H+��>�Bނ�����L�>�}���}��Lg�m�%���/�խ�m�Z�&���:�: �w1J�����9 ]��4�$���n!h-.��H;��C� )���t9���.���3�]�-��7���G�,W�K��0���^M����m7*
�r\a���qe&��wg#2Aq�*0@[b��*���HF�����o���mhk����=�n?Hա���F�R���o�,&%�&�$_�o� ��Ε�f�����,g�*H��u���7�w?S�+���J�?������9��J���(�C�0gw��ïW�>O��2K�p� סē�A��~�lJ�s�M��n�8!��E��9@L���u��r��B��tgs%fm�Al����ӾȐ�7���GY�Of$T�tJť��ḫ�����SM��a"�ȕ�G�ΝJ�@6��蠶�A;|����=nDֹ���]Ŏ�}P;3�J�W��AS<�I�QY����-�DU����`�VF����S
(o}T��D��z�t��� ���Ys�S_$�`�1��wB0�9�'�l:�.?��e�[N��y$�u��o�@~l"���1n�,�3 ���pe����t�p&��9�J���Lc�Rk��b�P߾�4���?���!R[㉳�7�����'�_f�-����(�٣+AaP���ǁ�l����e8dt�����%�"�	=����=�D�:���1�h�(��)�!�<����wu����~el�rK�A�63�U'4�?:���h� =��շ뺲��;!�W�B�es��Y��μ�v�� �.�3lf�F������ϳ���T�^�O�HX�'�_.�1(�~�ow4_>��5�m�����M��wm�_:Bt��0r'2��B~��+�<P�e�j�v��I\ݭ/V0`�۬��Ĭqѥ� ���3�)?��Gvǽػ@5l׷y=���dx��~�,�+gC�m�\[0pU���]�UI`����@e��~*ځSW�C�� 3zzjC  #R��1!�0!������n'�6�|T��f�H��.r/�q��֢U,d�W���4�dv�F���[]'�rN ka�A_l[�qY�;�ՙ���A�s�t ˨'d��ퟎ�5��k�AJ�NϮb	�c�[�T����Γ۳c��! ��xc�(��A-)�F�F=��x��e�����3�!^T��_�=q��C���s��f��I���>��Ϋ���ʾ-�η�ÿ���*�m.����АО��\���'�-��`#E.��|Lg9_�f�U�>鲢gU�>g�o��	w�7��\������i$7��h�ӭ
�9I���u���O6�;�d	J:�C�!�x�m�5P8<�Ҋ�{sc���y���9�x=~sv֗�f<������/so1��ccQ�T���e\&]���b�|���W&"myu��0,�C�q�F|���f-ٝ����.B\N�W�n��fD<59���q��e(y��{���qKS���F�V�Y��$�q?Xceo�ߤ;��9U8��sZ"豴׮e�Z�'d�@��kU��"�[����{�k�-������&���u2ض�*����|-�K���8�[my�dPQ�aN=�3���0�z�������`��"�?���޽�5M�^wmg�ӷ]/�Ȃ�LV�:a:o3�y]����7��b�������[�]��'�����Y����w���-�|8./����8��Z��ϧ~|�\^��p�X��;�a���x�{g��'�	�^3K�hMط,�5/(���c"r@��Lp��;�c�r����&X��,�Ŕ��YFp��iI�;6l�[R1�L�A�)����dA�0�����]�dt1���;�oݨ�X��.�/�p���>���THK:�Sntm�"&*���d�@L2���>)5���SQ����� F�/B����P*�ޱ��HN��_�Z*Y�<s�k��!�"N���H�	�=e����naH-t�X>t(t
�j�M�A��߻p��,�F�%-ٗ����(��8{��I������I��D/ sn�E
ۣ��]7�n�n�q�'.1�7���?+����M�f%z�&M�9��U���aű$ht�|�k���/bB��zI�K�v��T�G����?������8ߘ\�<�y�Wx]P=��1���?��^t8Ȃ],(��&BH�3wǯM�Ǎ�>���:s��%�Yk*l�3D6^�!����45��v��	����1h�Ɋ69�TɑaD�,deL� �D���7���Ȗ��@�����:mL��<v~";�����-$�ce�i��RK���'O�-���[��-JX�%���U��x{G߽���&1�������`**� ��;]�&m|X
�e2>\�r�[[����W?�\�]&�T�?ą ��q͝{����2nk�Bu�.Fo�O�B(3��J�D�U�I
\!$�׋�/�ް��'=��t������G]��WP���m�H��
=��ж�Z7�����h��%�C
�?R�5'��!O�/���[�س�?cѨ�H�� �o��Ӫ�D���Q�-P!���e
�[b���-w���*��>��v��#�OrȌ�9gp��}��|'�!���� q���������\�w�Z���;#�MFl����}*`��BK��"�O��ΰٙ�ajZu��f M�n������ǵ��V�o`7�hX��)�L'4j�k��h��)k���xc��~�V�"k�����U���oH��-��r��!��A��<�P�'E���+�������i'��z��m}��7)�t�J�Yӫ�W)��ǀ
��񊴐�E%�\�4c��`F�����S�yUL`-����?ճ]��C"<Rd���,��4�I�L���ɲ������1�}noL�&'��Ok%���YAZ^�2��u�Ҹ����g/���7����Khr�v��oʙ��`�YK���))���a�/Ai���y$������rv�迥X�vW����b;]��}���|ޏ�..LCF
�`�;B>�Г���%������9�X3%�'�����BjȎc�m�WlP����xe�JV�l��߇�z��.2��TW>a��a�2i.$:'���e��rh'-�����;��A��~>��R��[���)�#����J��d���z�>)�\6�45�|��",�d��8�2d�{����4cNk:�*�{�u��p��A�볥�O!}a�`�/\T�h���K�V7���&@G�妋07U�!�$G�Ä����q�Zo�#���
a�\C���n�*������5
I}�^>C��|�֭�a*&~��-Z�nL�L-�� lt�ߣ6&ϸB�+r���XL�������w����cGL�Bz�j�,MI0/��4WW;���O����FK�$�Q7A�%E���r@�+Ԓ~[�k�jF��IB�`�+˰k��V0-<�g�g�+Ի� ��w�*d)n��=ZQ�']|LL/Ip��7��>�6@������=�s�a���,7�@����RH�e�t�S2���ef�+?ܟk��AK���"�n�O�5k����������*m�)[�����'Ϫ{�g�I�*a0��E�̊4�W��j��ހ.F���{\u��@��Xm� ���Br�P�C�.�x�~�$�#^M������U�K��`bj�m�ް]<�]�.=�Hٶ�X��h���5�#�4(��vO$t�y��Q�"�B�TQS����?��ZO��Y����$5��O7���č��N^2�S~��������B+D2�����D{����w��WA;��%q�l�}}q?�hG���usb��.���P�x�^�M����xR:y�@������'���+�{�#g�:�(�ř2��'h�a�/E�;�����Z�JB�p�x+9H�6��`���� �}~�����8�3��N�r��i�%��I��B׿_l��!t�Kz��S)�9/���źN3���W��p���x��_���R���x]����%'�)��b�S�.�W�y�T��!?FL�1�`w=�J��p���i����z����O����bX�S�u�\�`z$�a�b��C5�K�����[F�,]Ã�������=hpw$XpN Xpww����������?�:����v��]=m��R���nI��/�d$���PǞ��6� b�덜�*Ib���(�v�����*'C��B��Z�1��R%?��J�ǀ�� �Ϛ���𦶠�����ޯ1�8�J����G#���k��4�[���n	\�e-ЭE�#yZ+.��̞Z#,���@R �#v\D��� �	�3�Vm���R>c����H��l��on�J�'���[#�y�A�ᢄ�2{3�
!y�P���G�LĈJ��}ʔ��Q`��Q?|�������.|�oɔ��߹�mr�2��zlT.$��`�������;c��3��W�#�:����-#�	^�@d;�'_����Tt�[���ۥ7z�%QS0�J֛k:f�N�s��v�^��#�%���?1�m���d�fO�;�p�f�d�p��fZ�FS�AܱcЌ�>E����r �j��M5��gc#��%��wzٝQ��l�k�u�m����3�ɸ��3_<�v������l	��st�wS�+̏�V�f_��M���1圜�%�ٛ���o�\�tnt��R<z����W1��w�e8�:H.���*Xs�{������fw=�>�[�k��u�'�E��J�4�1��t�8�S0�G`�=�x����nہ�k:�Fa8�	-b��g��W���	d5E��=� B�T<v6>SV��������$���8O�8{/*����$Fd�h�f����Y���ꝫ��D��6M������x~��k�%���F���_]��d�+��5�o]D�I��B�R�6�<��u>~�T�����Y���-f���Oe�M��2�Y����#~|_v�}�+e�-s�UN�C��A �鈌�D;nN�����j6���� QWCJ���n��E�ߙ�59�}��]�힜�_�������0�۴nf���L*��I��ſ��!y�W˪�b]���w"��S�ؗ��������o'g�`s<���N��l�qb�eҊ��#�W���K.R�דy�gdy~����؛���H�C7@.���o
JJt��bN�[b�?�	s� #/��]�p���gW�x/�`tFy꼝����������'cVc��~�Ww�f�U[A(�V� g!�\��ʹ`��-����]�Nכy	�����U9�`�4���s������[�w6L��������vX�&|��Q�΀���՚�b5�lJ6��˶������(��N��19�n���?F���ӿ\�/0	��h��U�m^O�CA�XJ/]NP4�,'^Կ���U2�͆�Y�B����g�y�<�K1���|Ϫ��/�rM��q_P-�����C��"l��`���U�p<�"� ����R�ۛ'&&�OoG֌�E�S ���_���qZ@�~`Ǉ��I��P��r�~����2����]NM�A�m��z�+1`'������G\�G\�k�:�~3���S[g�;(xrZ��y�z�z�ƗR��xee�b�v�1L.�%� ��Pu��]���SK�AH
�3)''ʁ3ҙ���L���[��~��|m��`i��kZ?�oe�����{1��:K��5NL�Y������^���]��:�9���S�g�y|t��F�1�%l~'d�$d� l� vBxǣm�MH.0>"��l�G?}�t3C��-tc�ﾧy��1�k=�ն�WE��u1o�����~`lw����:O��)fm���3'OȠ�j)l�!��z�gd�����)Q�R�绗��`-/�'|�SW�O���;]�}-Cl�.��f���������5.���F�L+γ�1�AF�B5������/�릫U5#���hI*-�����5�;�b��E��A֬����=�-�S�*T�޴0D9G~a7G�B@�um��v��� O�8���ٗ�"�#�AZ�!��w�e���5�"�F��5#�VP{�z��qoQ�.�+��t����]#Ԅ\>��x9�[K�S�G-��-3Y�W>�7��|���0�Z{��F��6V6�#�pn/�|�W+��?ؽ�M��ћ�u5��h����&���ր�8~]�Q�ύs���#�(��|�R����l�e���5�'nB}�{�\��!9t)~T�]�����)�����TW_�u�h|my"lns�E���,��S� b���2��(jvD#�������o��׊��^Y�!�<ҒO�Ee������#��l-�mh�or��9��������s��h�%�Nc�L�}�Ȏ�f,"vy�hjR�`�N�0=�dLV�)^�t��3"~�c���:Ä�� e�d>�vV4ߋ��Wȱ��Wn'��/��UcH;���g�B4���͛b<%�����@���h��2�A��_P`oV7A�����i��*#)��g�N�o9�ʣaT1sEOy�M�u���Atoe���jħ�vX|���U����X^���]�m1���$����A�.T��ԙ�'���� �K*�\ĵe,Pd,@'+2��S�k��F|Sr���C>�9�W$"�WRBu��L��	�g�A��_�, �B���Q�kx
׍�߯�ս\J��:��[4=��U�j�`@i8M�����^�D;!	
��}xO�o�Aپ�-���u
#ᳱaI�ʓ��!m�x�֫MA�QS�dQ'���ʴ��2��69�P~�cU\#!؟x��ۮz(�)��F��kӽ�o�߫��ik�D�dS=ї�
�m%��&=u���PL�Ծ�521YY+{�������-6"��O#�GG�����/�LmYɌ��� �E�Mx՞��f�-�)�|ĳ�;���"�w�R��t��W4qH�.��8 �l^^?��������͓$3h��_�i�Ah$9����%N���%8��d�Uّ���AD��*۟?"�YW��UIF�Dj1%%\�%cd��9R��N���o���;��Y4��7׿˰8Yаd(�� ��o{�
������.��e�@���Ō5'�hJ���d�im]���Sag��kZ�^A�33VSQ�e�)d�f��=��(&��L�<z�2�Aj?Z$�+��$S�dlѻ�N�K�|qHy	�w�/q����1´z^��q���d�O���(ؗS���B�������,e/H�P�}H�I��<�^�)��A�{V��>@^/��T��� �w�E����ܣ�Kz���XV(��}�؅8�cLv�M.����2��F���G��,.�[t��bcK-���h�ⴔMe����d��O�e_4{I���?���l�ުW͙���u �F�6�I��ǌ��m�!���=t�`%��\zԳ�FBm�lz�Ln�S�.�U��ԕ[*�_�#P5��S����U�TX�%�[��~�㣟r�;*Q�.�h��ݒ�i	`��F\ &�߇:�Pء�>"@Θ�d4ЀZ�t����gg�as��E�,m���?�>�*��3�j�{.�u�ph,1f6����R�'�s���d@�h�'Jp��ښ�*����@,�N5,V�	~��`(��O��Z�m��QK��L��j�KĒ���X�r��oV{=��ֆJ���W�2 �ўa:A��o}20E~ak�Vᴍ��Z�Ҳ0��d�S@�\��J����q�&&n�U���*Dl:��K�t���`�\�E�wE�r���WB}rɡO6���������6s��g,�ԙK�@��&Y^a̼2���޽�Z�*f�~��u6���i��ԧf�|$��t܉;����2;���?H O
�@Њ�y�M�GP�6ӔJ/c�}`��,)B�I���i�݆` C���E���A� U+.�ʕx���ҧ�˕so���d3�=��H���g�@�cX�lN�L�|�n!�L.��>��?o	��o.�R��@���$����/^@/�Q��˰P3��k�T��?�ǹ�Ͷ
��rI*�GK��������J8p�P��[3D|�������y���/_˒�Q��T�L��Zr�O[(_X�Ͻ�h�^�e3��4��8L]"݀i7��!���‼�¿������Xܿ��!��O�w	T;{�M&-�bt�8��7]�ʭ��	���Q�~�!�b��b>�s��&=3��{�T�����+KsܲZ=jL%�D4-��X@���[+t׾N���in�"C&t�Ǹ�^w�]f�����e_��:(*w����6O�P�e9�7�����+��L��b�(�mĖ�����?Ι�I��������x�vlff0ϔ�TZ0�S���>����Ң鿫hݺ��#m�Akhߨ��흽��
o�wϗ�Y����%׉U�T�V��|Ig}�8v&�|��L�q��U���3���5�W��m�-p���n�ħ1�W�;6��,X)���LE$(8�!�2�-���VP�H����F���o,��e�Vi������T(�l�ڨ��3��l���?�4�ٞ����F'+ʶz!�}�ne5l�ס��z�Ұ���y����n��eW���{�{΢���)r��.�uQ���!;߷S�i�`�B�l:�d�S_�m.T�:ۏ��8�7;��e<��b)�kp��D��:�Һ=�H[�{H��RU�N����~�Z~=��-0�?�s�z���Vc��M�ϗs�U��/����L�9Ev��~CP�X��n)d�j�>M�
��U�q2L���� �=�3~�W�C��s����M��ҶH����6����J��L��魗�^�ˏ��|�򑢚s���,���~���Fa9t,�|D�=��8/3ª9w�.kxT�[c������a8ѽ�Û�ն;׍ԛU�����J7I�c�sJ����ޓk����z )��$>�|B��¼�ȶL�N�Y[��z�f���.��c�yH!:Ņ^>�t2�DOrO�	1���!u�����j�#��Q���%X&>{^=&>�(�֠��b�?�Y��e�{)'�:�5p��[+�)ƿķ^=��Ԩ��~Y�B��wЃ�c��zk)8�7CjT��ኴ4��Q�����PZs��ع��Y�5��������u���*�'�r����k�;�ƺ�^��b��]�K~�_�xH<��=�K��B�H����K������y�o�RY��|_8��
&D_�6�6n �/��_u�徣É��i��l܉oڿ�NL�p"��\�q��׮|�������۫5��'�Z��I���`�{B[��Ids`BTf��& �|a��Vz5!��jdJ����~zE���DZY�i��0�fT�NK{���bo �"Y��	�����3�r|Oߞ�F���ڷiB]�P����K�݂�s�~S�+w�e�Y!M��o`�U�_;.��t0�n��n��{<n�~�����OY��J�=�0��� �����������}e��E;�d̈�:�b
��gÕ���plJ)�N�����ߝ�_\�8�����2v���c韧�52�rӝ�o����|����	�u���B���/�=��
�@ �X�mS���R�f!sy�A%��M�ѫ �"�L4ǑԴ��Mc��3�������WRls�'KY -Oy�Y�i3�i?�~Ww�qB��1E�*(G�g̛�n�+�����z|�6!ľx_���{�π�s��0�wߖ���$���ɋbOX-��Z��S�v�]�w�Uc~�ډ�b�O����v��V[���7=�z8��:���b��
�1��ʥ�3���Y�Ғ{y�tUo_S�=�^��x�Rܓ�E��V���t��[(
f�� b�*��l�z���b���'Լ������ ���<djG*�$t��*�u�kr�����g d�� ���u!�l֨

]�L&>-Okχ'_�T7.����z�h�������o	X@�J��"Tg)/x&S���Ĕ���QN�θ?�K� )��}��k��-��Ѳ���&(ǉG��p'$H���3��:��_�U�/�$�E�(�������Sz\�G��O?ɷ^&t���|
w��%ū�W8s>�/�];��8n"q�ޤ���&�qh"A�6����DT�X;;�e"B�8_%-h�s'��ʏ	��É����c����H�d��s����^�&I�ѹ]ٝ�����e�-[m�q�M����-�
�����:tR��J�-O{9{�ө��.?�V�ϸ����'Q�q�����Ɋ{=y�^k�r�$}j%��A����ű��e-ؽh�i��y�|�qq��jY��H �۲x
6���ò��7�����J9X�����rȩVQ�GMX+�F�m'�5)���d �%/%d!G�z����ix��j7+P�E���Q47{��H�=	��B�N�ʗo����V�R���!�.鏤]B���<Z�̙)��g'ށ�e���b_.�)� ���~��[�xEשz���jӤ���}n�S��'�D���������*#��~ik�*He����e�Q\$m~��CzB���W*��ڗ�����kq���m\�ɳ�P��OQ�����|Q	Ũ��᫘:�n�4��i�i<�>�S���+�u�z�?y�>R���ԥ3�k�J���+<Z"��x�i�I�E2ђ���s�#L�Ղ0�˿�v�ޮ��}���+�����1��_�M���@{�B6:;w8�M��=ݻBtZA�J�r%T���J����`���Y �N� \�_�+=B�|:p�%<<��������E1�#n�2����p�v�;��P7������K�*H�i.�#簈:�ބQN��=}�*��hl'�r���S�����\�p��-���)+�q�ϛw��~?�ヱ&`-U �P����@5�/i56���qӫ���ul>@��V�RzR��R}����C�`@����� YP�#2�@w�*̅��3",r�W���ApϷ`G��f����X+u���|����U�c>�1�N����Y���(U��t����/��^r���J��\����9(�)�����vFif�L.��3�Qy�02���<���җH뮞<RIK=���֕�/)�4~��֪(���§��
�К�%y,�&���9��qP#���%����1�Y�t�V2�K�:�������0��Vyx��������e/Eڈ�1s�۳]A�J��	e�ķ˞�<ᴌt������`P��k�z��WU8�&���`v��7�T��@��Ć���k2��2�̏�w�WgQW�*��$�o#����]K ����[J�L�'ec�t~6��פ��JFDN�S����6r��u�M���)4}�dU�MMZs��4&�<-�y�jB�m���3L����c��H�PQ6}\|�r����E�Ŭ-Z���p�t�k�&�[5}��5��}�8`w���y�5�����&�`c�A�Ʊ7��Py?R������2%�:�/.d�Hd.2�s�_�=��76�5x�B�_���Ra�MN�iR��6����~ٯ:��,k�𽇃M�.�FNG�O�c4�+�($� ��Q�����|]~�9�WHh~~m�Q�;Fi�P		o�ҺX�C�;c�r�p�u@���>�}�z��h��Q	J'5ux"
�w1%qsa�?��ް�G��吘�ż�����lW��5��&����-Po��/��(P#b�����f�--e��ы��#�d4?�ֽD{T��Gr�s�^^)&���)���iQ�Ҽ�[�.�>��ʈd�v~��#n𩭻gzo���$5|���Ԁ�E!8/�n�qhs�]t����t����gc`�����Z��H�1:��˒���>�z�4횊p����Bf�zn���	���v��	��HF0^��^! �R` ���y������*�j�Mh{a�𩖧�8\��dlO������!}i���WG�]-Rw����~�����\�|j��a�O���>	�.g�Ռ1�����i�?�%7c�MzZU�o�6�e%0q��f^�����M�~�Wg�
\	؝���%��o��z���Ⱥ���g_����s7慆��5<��?�bz�������St���G��*���L`ڴ�Kce��O��V�d����.KYi��	�O���z��cߙ��5��OI* ��s�i���B'�(N;K���Io�\ek��T.YlPD�uM0��Q:z<&c���*�(�Ď�,b��1`���3@mQr�`���������~���5>A��B�d��\V��:�y%�r<��Ɉ
~>���Sh%C�jr�9K,�a������5i8�]zvs,1��\��z�B� �}L�P6H����*�/\�ŷ��;t1W�n�|-�Y�֦ԙ��j���ޕ�h�wx���8�f�$�0V��L���#�8Y�����IA0�L�\���c�3_�f�6����"�����C������y;R��	�4��0�H[A����CW�f����>��Co?\���E��Ĵ�7g
p�id��u\"`�@OTT4�;��B��/�Lu�h[|�$56)���ت���,�E�@������A�;b���G�9[�rd�I:��f�{��3����۪ ���X�֫:���:ƪ}:�����%)��;����Uwp��NDn��e�x b�&�o�p
r�J8^�s�Еe�g���8�&� �-����l��X�ҍ~:�3���BQU8�5·@cV	"�I�)�
1#�Cb,m��T	]�٭�g���}��z�ɲ�v�����*������䒷TO�{�y\_L��_�HE���Ay�]d����K����;���_%0z�*?Y�
t�9w]ꗃ��T�(N�慿���U5��%:�"�����cE��v��[��O��*�\���A@�Qܼ�t��?c<�?�Z!"���Ϡ@�T ��8Y�D�l�4���l��eQ��(8d�^��Cu0���7��2���u|��}A}ը�1�ر���fH��Q�ǼԬ��m$��N��7����wǋ�}~-�!!�'E�[$Q����\TcI�$F��c.�@����q�u9��L�G��C@i�՟� ���l+�����Z�v$.?c9"$)�Fe]���_=�Yi�V��g%|�+�As�UR�y�t�/����fW��=.j��kV�v���4��g��yc����H�X�Z�c�MbEg:^Z��t@��'"������l�����Tgw�!VS�����hW(#5�dBa	4 s�h��KO��n(��vL1��蠏��@+L2Ԫ�+!(�B�!EV�a�X���N���੐D�����;���G��w
~�6��+꠆P�Jܛ�ȋz�����W5�.Jġ���cJ2�!C,�,[?tG����fW�{ɐ3�{��xI�y���+����׈�޵,>�$���@c^�M[������)6	6�@��ܥ�����x"`��m���M�5�m$��͛u���8��� ����W�j�z
���v�~U~� ,nN8P Ԅ�]3���h�J�����6���,ץj�x��n&�	��;���� 	j�ٜB�� �V,�$l�G�<B�qܽ�Оj�[��M/��!C@��	𱧁]�_�Y|�3��r�k-�!�]�̤g�~�ط-g���--x�dR�u�e�2{�P��Ix�C돒���d�;uʌϛ�ס��'��{�F�������a�$(����'�"F��Y�0	Wc�:�8.G��*�C������&�1x�p��4\��lbP!�G�c''�]��c=J��Ve�4�蠗�5M֕���p�6T�ax]�B�s��IL{��d|�󃆉�-���#��[JA�(�>�g}��CM��� hS0:����[lpk<�{��Ƹ��A�mbJe��`/���UT�\+mC���9��S�'���e�������<�����f�)_��[�e\VUM���r%8����K�s{�L
	�I<?��J���^�{.2q�'��M�.��, L
ڝ��E�T\Ο�qqhFI��@1]m�*郲�/��|�?�7�I��f�T�p����E����C�P��3���Ԉ�rb���6�S���<ǁ4|�P�:���HJ�$D�S���?H!ㄱ���WN&��#�x®����{]�b�G��h�D�hZ�tY0.�ew	�G����h5D���c_+IqR�t��TM����ϲ��(�[ը�}'�����}���C�ɉ?�"���a�u�%-xu3�J���>�͖[��z@�Ȧp4�b�'�vQ���z�����ȫ]OI�����r{���x(������M|��p�ts��f�LE��D%ASj��ĉ�-��xm@[�WṭjXC�%j�\93��Q�	O�i�.� ��|���KO��?؀V��n��S��kz�Q-��JǴ�g�����sM�ͽ��2T%�'��%V�-6v,G�(�:�$�l����:�25Я���V���ڌ	�>�%�	'��h)|>{�N�M
�ّ���P��l��&h�Z��Z~�}o���C���b#��.��Y�o{�7m3�9��37<������y��R�ԟ���s�74�UUd���E��r9���?��n`U��L�)E5OS=�_�(�o�b�r��hn})�����F��A����B�R:p3r��{��v�����g�W�t�c3}"=�WgB3}v�?����l������܆dY� D�%4������B�H�x��%Rs����8�>�NXmU9��ן/��tT��ƒ��>��I]�cC�ӈ� �ƚ�U-g�=4O�m��hN��pj�s☠��i�k��r���%N�Y�|y[�7�kD�
?&$7	�r���;���$foq�h��d��↭(���/��@%Ө��^
�勒�����aJ4R��4��=�_����w;����)���Rb0���z�}�8�y��]�3�E���Ýlt;�ʄH��4�I���J��n��l���~%X@k�ꏷ(
3	5&�_r�aU	���EA�U�_c��H��߸ID۬|��$�a}�
/&�([|5ъ�T;�^%������o���e�U�x�h�����Opg��m��w����=wzK�f���מ�;&���3T'���h��o�=�>���'z�@Opn�Z�yU0����n�E��Ix�w�k4%��&���|��}�n�%z�U��6l J.۶h��'�}m�,��=���G��c�{M-DE�%}�L��!O;0p��(�(��!S�<�̋�$��|i������(�`R4�r��	k�7��η%H���7��y�K���I�\�����xm'�I�u�si�M�QB�m��rg-Y(t����r�s5sBE�ge׸ǨJ����Lfq)y�B��Ot��u�6O%`,=�ׁ��EP�dqԁ�»�r�t�u;��1����d��b�/'������S�h4-����|�[�^��	75�0XO�x<� ��<�g�D�>5�[O���G��p�j�:���?��7�����u=�e���@���IF%�a��"�,b��9�b4���;o�����}^ŀ�av�ߔ��G8�?�7�b�y�	�+�oB�Cĵ�}Y�i�?Sbv�#+:�P��r���t� 2GG�����N�c��CWU:�g?u�8�#"�>���=Nl��K�$����sb��b�e'��
�9����2ji1�q�'�\3������'�M���i�О``��Ɠc]�}�@��cL��U�3��<
�2��c�����9�z���%,�R��_a��2c��kkf�S�}�Z��pm
QV-O��MQ����9��/���|\5ILֵ����çN+K�x�_�sɫ�R�<�s�X���k�&�S:i'��܉��;bObNl�&į��-��Ʉ�*j\V5�i6�"�����<l��Ծy�gAI6��T�]��^����/,���k�[A�r����9&�����}��o1��D���C>"�키Iv���.7ԶM���x�8a��Y��}`>&��?�;NMi�q�4��[�B5���ߒ����B���4S�Fz��#������0M�N�l�[/{�(�g��O"�8Ԟ����2C6ʫA�����q�ۯ�KaO��v�ק�#*'øXE�X���X���������:��Q�Z���������v�HJ�\��o�K*�ej�ncu
r����ˌ[��U[�i�N �R?&%�����DAAD86F��P�,g��G:�\Xn!Rɰ�*�"O#kq�;��E��>]�w����+��,m�P�tG��)T62�)ahSb=l/~C﹗L�#<�G�>Z���/01]X�ͤyB_�y�f��`J�\�x��p1�O�Ard�'��2��_�k8n�W�����6V�"L��BǇ������y.�ʋp��ݰ��|�
(�|��Ib%JV�~�ܻ�t���EM��|��lφ'��:ػלg��$l�"l�)B�&B�G�^I�LI��c �.��
�a��)�n�	��E��$�@��GU���铫 c: @!S�x�� �&�����d���@q!�����Ju
<UA�5�Cl�(����I���hȆ)��~	�
-���@-f��s���G�#�V('�O)Y�?��?�_٫^�U��:�_���P@IT<�C�Z���vp���+! U�זvP���Ό�t�ދuN���L`�w^o��Xxz������VPLD����X[���24�?�z�O.���{B»ſ㟑����AcPԻA45BA���`�x����Ո*^���]�9���.�Y/'��f,QnT%�e���k�\�����w//�$m���_��P���)�}t�l�1yx�i<�~��W��)��\o���<w{�3;� A��OosY3�TB0&O��{B*6�o����($Ԝ�r+ ��,�O�!�>\%�H����������ɘő��c�@�ޛ|3��x$�s�����}��I?0v���t��*>�rT7�A�d{��
���=<h�B�q�(^�fGz�W>��^�� Ӗ�U��p�����������
t h��9�Y��R2��2b�\I�K�HH�*I�ƚ!�g��JZh轾��@9��%$� �$��1�Fw�F�!��n� �\�X2���;8�S�����(�c�F�Yԟ#ɱ��=������6hF�i,�����Nޚ/��R��s��� �:��*����dн����h�t�d�47��_=:�aUqC�k�X�k���c"3��vP� ���y�,�f
c�4�.�	&h`s��0�����Ȅx`�@�3x{���aEM�T��A#�ؔx8�&!�\�U����i�<����"R���y�04�"��P��Լ�rj����|-��K��`�AN=	J��
R*��xfk��P�|u��^p���E"#7#��qt�G�j�4jMZ8=Bh���e����]ӧ�d�t���@����f4��[���3)�)%�m�W�)������Z�m��SY���J!-,j�j0�{��!,^y��(%��Mh���t����W��l-��M�t"{��a�
G^Md|Sv��y��F�t$�$ªؓ��O߉/o��T�Im���߹����7a�y_x�	�
�`�[vG3�C�6����	`^�����o�?�A ���/[K{�m���;q$�)~F��7�l��R���p��r��e�Z�m,!T��{nѾ�_�9��E�3#_��5a����KЭ��\�������Q��e��(yd��z��m{�q9����Ø���4琔?�p��F�Өc�IF�)2M�M�u�f�Γ$���8�V�Ӗ)`� �/]�|P����*�Nx�Q��܇f �m�1�Q�{d^�VK¥���N=�d�aNF�^�1�\�ܴ4}�t���S-��D��$�OA�G#��5���{`҇���'P-�1ϰ~��g�`:,�}��� ��/�M�.��VԼ�I��'��J����=1C�;���%h�f��m�P�*���	�@}.�6��&�-��b���ɑ����z��tp�a���d9섳�$���
�h
���"�讽��a�mZq��(��ň �)[.�X=9p-Th]���E%���J~_n�VVs�7B�KU������錞��� ���o<��l�m@F�J�M���_��}q
�y���W��g�1�}�Lb��/���\W���No�}���m��eq���!�$�1��!��s������o߅�nC�L/��,ω��>�>���v��=�oÄ���p.��>ȕ�(G~ ��C�\�BF>G�:�;(N�,̋tۑ�vz:�hmZ�#��}����X!(y)���{��$���`2�`g�g���-u��lh�i��9d	�Ӫr��|q��݊���gS��(��عq��V���>�v�Y���<�ޢ��8'�"�X���2�o�Eͤ��wJ�%6��GV�烦Э]o~���o���������CcL�pN�a�ݒ�7F�p�c@��:B���V7N���+�>�ݟ0���f�L�	l�_-��k���f�?Y���雞�h�\�G�(�q*��{�Z��*���JH�g�p81�p�F>���¸L0+�߅m��p���� �֮��<NB*	B�"!�NA��6����E<^7�:0�h�o0��y��a�ʉ�Į:���UmT�m>�Q|s�c>��n��1e-�����gf��t�˷��5t4��ު\e����Ɔ|���#.w�Z���x�����&| �J:���b�|������n���6Yt��;�2$i)5�Q����"Թ�a7�/(移��r��b���L����8P���:�t�6m�d��7׽c$�`SA=i����>�e��>{ �D�0
:���z�MG���#��1��uy�,�e�2���6�. ���Od��=�<�)Yҕ�^prhm7Q�m���|��)^�I���\&��S��c+��@��,�-+��#��\�)s���pvo5�~>!�ݭH�(8l��#�z���!qɧ_�{�w���-�>��S�>! ��W@k���s-)���f��?�̧m�!�E��"�xY�&�T{(�T��5��(�0�k�Ow��ΆPo1V�����e���^���b ��+����~�R�wuXY:�>df����;I	��t�	�D�h�`�X9P.�̞2E�3���"�������$ c	��ٵ\�>3մPK��#����]�.�nX��B����jN���R0KY��|P�!������q��O�ioB>�t�lX+�Pw��q~�=��Qz�E?NV{��L�x`x8Nϡ3ў�<ॶ�e?0�q�f�i��F_�A �i�9�(��?�y�11&"��ڂx9w�mC�+ɻ��
 ������o����� ��H��A����p��z�K��������:�24u��a�P^	�Om�`�&W�h'�!��O�y `��3��=�	����Y+b����i�a�X��t>��~�, rV�8�\{d�9����;ٵ,#���Cn�v��vv��\�E;�Ч1�׫K<�_WԱ ��C�	z����6��s� p�/+�-�J��!O���`M�����E����M4ӞCl�Y���kL���+�._��m֡����:��;n��2�5T��n^./=�y��ƾ�/�_��0�*�s����D
�4&Q��{��ϙNçv�>v�֩_��F�����O;����md��?qq[�C������Jz·���@��v�y|��0~L�y��>�|����3�!��>�<}�c����wL���V���Jr�0���Ryg��51�,r`lwX�RS�S�= ͙m�E6{TH�w�6�1Li�+�Y��4S��V%Gt�bu^yi{X@�A�
]h�%x���������)�ė(�x/h�w��������!�َcu��7��M��\x��|L�*&�����9�l^���؟���R�k�t[c�<�e� 28��}��~�׈�O?���43X^C��<1�����[]�RPP�ٮ�ڄ��Eb���*2$���bp�� �_���Zcu�2�Ͳ�r�`^n~O��`+%�b�1�0V�̈!�GK%o[�DA�\�������7��>�'S�Bs��3a����ʺ<QQZ��&��	�L�Hť��� 7\ʽn���jU5���Ei�|)w��E���ۯ�[)a$Or�	.�UI�����}��\�po?i��^�`�X�DT�"͌7��;��=ئ$g���/Hd)�B_�{<����ӕ���ʗ�7�8��G�1	x�7� g����f/(�*H�~���b��U`����g�}%h�R^k��2(;f�ݪ����#�43�T�R���hܟ��W5`��
gmK�5A�B�n�'��m�D��;�x6=qj�#���
|L&�؟[Q��ُ06^���N���!Ex>癁�k`z�((��L��'E���̹�ēȦz*���fWGM=��i��$�*�ST�)�bڐ��G�:����m�����;Gd�<ܭU:�WED?�N�wu[�d*uP��%���_!�lq0B���RR�f��Xo�H���� ��y����}qwwww�]����	��!��Bp.�'���w���W�UKQ5�5��}����M0r棽w����<� ^��9���t�>��m�����(P
;	��M �CI�V�|���s��[��	7��a�����װ�U~�T�ꋱi�
1�$�A|v����D�z��u��<�	�\�&ĹfՉ�<�g�'�i�{h!���s�`̮������f3~��w��v���I0;qz�.o{)}ޣ�;)����M��J;*dŞ���{���;�Y�:07X�����n0�N/���[]:��+��E#���D 	O���d�g9R��P�pxY�O�K
)x��F��1(l͊5����3���V2
�
��r��S�G�=I7�\ A���Z�3��ΊR�C�0��vz��H��+損�AO�kjfGUɉ���1�����ߣ����u��a��l��֐�N��Mt?���(��̪��y��\K�O�{�7��[@�I������݀�Aw�1�pWa�8�]�b�i;O؏y�ʸ�o���.� ZUj�����Tt`q/�o��޴�$R��l(G2|�~kg����aw��+�����aKρ��ܩ��33�_�G�@��Z�1���8S���	��p3�W�#Q����TDWv�iz����Z�;~*�}`��rQ�} U�wݘz:������hq�ِ�(�
�5��A ��
>�����!��',`J�r�J�)?r��Ĳ�#��0�+9+r`��Wo�{��CYߑ|[�Ml۱���<2��+]�����*v�`a�d�T������]�:T4��*�+Ԅql��VHɯ�9	�'��NYWqމa��D_�(>n��i=�IJ2b��$ڂx�sHU4��	���=����u1���"%�φIp�ת�<��nrY�'��t�m긯�x�b��0ط;����fS��=��~/��̅7��p����DD�ͩ�3�Zd��Ţ\�`Bx�����}RE��k䶺i=���e}�q��ek����=�V-/m� �'p�EƠI��?dm�jTl�� OnaU 0Xj�f��QQ`=9��c�vs,©Lչ���������
z��xJ�J��9���	 �Ѱ��A�o�򸑫�@��I�1�I��=������>�DL���v��^�&ʣB�tJR}??��$vр�q[�d���� yhhs����Qh1J��`0oX�)k�qK���Y����� �8!�,��.�8j�u0��V�fvW��S�T �EÀ�ы�ͭ�YB<���*p^�_At0��Aex�I�|�^��V������Qg'l�%�/L�w��w��V��D׾��ť�R7w7�Ad�����%,��d�Ӻ#	��o m�˭���M7��	.��q֖�l!&rZ�6s�`���Ћ[�4����a&@}t���mZ�iʧ�o�1���*�g�~' �]���tj\����xc�~���2?�������<��j]	�t��6��u$vsC{��Rc��q���z��zw�,,���_��֗4m"��#�j���5����@>�����ʟ�x�_G�(� 8�ļ�лG]�b(�P0�a���1��ܾ �J�( 3�|#��_���t~�<Z]�A��7�^������b(�6zngf��u���h>�t��~�W�(L)�0
ٵXWU���T�+�㰛 �]�fӥ(��1�3L�������D��[ޔ�P.�!���aLά�֜?�+s�1@��ymm����-Е^�)���'l�)���d���qh�Úx=85���XJ�Ӡ�7�fP���5 #����>/S���vm�?���{�ht����4
 qݬ\*�g"Ш�)�F�*3�EF�ta��� i�	?6�C� ~O�~*�B����C���w���/��H��JG+*[����9��H�S�af�&f&��'���9wKt��@�I^r�U� v d�?J�Xe�JqQFț�Y���Щ���zHmGQB��w�ܨR��u�;nЇ�qh���a�\�T��˅�������^+l�N�,7è�������e}�A}�D�Q�V�����m�*�g�@��b�����7���aȻ��;�?�8�n��$v���k7�����o�î����W�=��4
9�T�,��y�i�@��f}N]�?�\�h�d���k��16����0E
	�e6_����\)p��Cc�x�3 ��j����D�DE�Dn���<�;�bd�ڻ�h34�8]{�+���Q��x�W�I�13	#.շ�����b����j��-K�uU�w�Oڹ�U
^~�å����K>�Qd���-� ��[��_^��}W>�$E��ap�G�R�d���T.���H�,��t8H���R"��|+��)�ϐ�5�;c�Y0��56�\>���"���#�������6���o�XP�ΖdXA�  �fU���N!=�����=������΍��!ꇹ�rghp��uuYm\T�>�;������:vշ��v�h��G��!C�r�.����R: )�����Egi�Wn[�)SR:!S��jp@�լ���;���>9|�&9�t���v��ҝ�[�rXB��"`#�������"�x��7�:!��k�¬�R�������9����H�h��QF����3��M�t:7�bv%r�.7мܾR긾3�ߤ�]��1|�FK#��%,�?#j���{?d�QM��e=~��@Seƪ&�1��dl����V���y㡖A?�ğ]����
��C�������0�a���[����}ƓO����?��n����K�u��+�J&����F��������Xlt={�S �.�e�ٲ���z�F(�xϒ��		H-Z|��sy`�����ܽa#����8�A�bTS,pd6�x_�$��l�Ɓ=
;�o���ԟ1?�V �~�U	��j�v2�a�)��-}�'nU��r��USK�y�C��N�� ���>rGώ�m���Nx�$���KD��4{R�"<���Od��`d8VI|��W��M���v:�Y���n�.`?O7v0��p�n߽<��P�43��F��+�W> 4�,�*G�ӣd��6\�{��;:�1��d��쿦�z�#@b�6����J� ���K-{�����M:�A:<w�r"㌛~O^~�}�!�䜏Ҹ�\����`�bDt��o�����)(%��(<9�a%�;W���02�7�ǜW
p��^MDk��|J����e��ݼ<�H�D�q�Aaa���߂��{k�C=\آ*����Dе`�DH �J����q(2o̴�9�0"P�S����{��n���Z�z��3,��Rkl�/�����2),�M��ֵ7��2_� �G`[���J�Qa�����(@)��JB��Uy��������W�z�����åu��q��Po��睍��rvN��}}��ã��C& ���-Af�H��tr���O��v����=�}>թ����;]R��t|ZY�"Ȅ\�d������?;Yb�c�Il��>���0���>ƨ[^���r��25>��]���?XM��-�S��~����sXf������&f�+���_�<��40}:N���}����Bå	/����}����K��A���oh��wn�5�Ya�3ɑ���më+1]���>�X>�"�0�лc�d�,�	SSP�y�������Y�L����X홓|v0��|i(�� �>b�g�W�ȋ��^�m3%R��I�B#�FIB��PR�YH&*sڝ�'n�	ݑ�9>�*s<̂F@�Lq�y�$��~p�uR�]f�`�6����_!����d	���}�{==�6n����}��r_D��n��NmHꮇ�z�fCn	��y���-L��T&�Wbb񚬽��
k��fq[6��46���#��!���T�������@"�`�� �� ,��6�\���	aL\�������B���5������~e7$K�K\"�Z��n\�̗Eڊ]\?k�[�I�2�y)J�4e�X7����=�����Y9��\�3E�͂��W�|��{�n��j\	Q����)LW����D-�L�E!��!T�F� g7��]��O��c�a����]g8<�JB�b����O�����Nṇ`L+��˗�HƢZ��a\����\BAr,�����"Dy�ZÇ?,����3n
&�g<�k£��A�{✹EƠ���s�74v��D*��ړM�lᅫȡ'������Sp ??�|�w�̀I�T1ds�r�a����� Z~��*�<�p� ��sx=�.
9�}~ Om$��"��"�$wv!s�h�A�r�W�7���|E��Îl>ey%n�2�2�9$��H3����ˆE�_�>��?N�i��N̈́�
�z'�>�H�䀘!*y~X��T� g�i�W�$���{}�@n1�T�XY�R��&�ۏ&���n�hD�� 1�e���c�
���M�ġ{��\L"!��� �����ņc��h�AY�d&A��[����ކ%�S��c%�蒰����NU�{h ���y�����7Ѡ��x�"P��=��8��?V�RA5��(���N�P���)�B
��v��w��U�7� a:�`�ì��ހ��~\���:ðax�V��!B�c��w�I�����FU��?[��*r./tL���42@^�7���8�����~Z^VA���3�A�Ie{
8�V25�*/oZ1p��}��;��6[�����	Y�����Y� ����Gb��L�#I�t'e/9��/��ގ�q;�胼d!�bN�K�2�̚F���c�F���f�v�w�ө�[�D{/M��4��Y�����X: '�����R82�_����u������ϊ�5OV�
x���r��ת���z̬ɭ�0bm�Y%��W�\���g���B	67�y�Z�r�8���2�O�����N,!�7�ukh�>�d�f��5V�8DM$���aÝ���haa���C�M�hav���w��ֺu�R#���i�Y4�=Ɏ�/���?��XFnor�x��r���l<�Ή��|�M����MɋB�<�?>���8��D̳�k;� ��vR�!���p=�+0F����`��X$����L���ӈJ��ۙ�0m�Xj�>o�?<�A� �EuP�v,�d����ԙurqK��I6RcpE��ܐ��]�Hz�Q�+f�]��q�>�<����#w��w��L�s45v���&�IMO�hmV���gG^��������wx1�Վb�E���0��D�,��Ww���-�5��/7&����-?LR�XF��(�i7sV{ArP��b?�,ݬ},72�y<P�Ӆ�6G5Y1��=[Q�	��+x)h�B��MuҰ͌��{�<��W�q(���	uRc��IU�� q�%���^�#?��龀�~jVIʊ�� l`��Š�1�F��ꊞ���AV8��ږ G�E��I��1����B�&����҈/��ǅ?!�w��lE�����ɓ8 ����'p{����d�yh��Ï{B�l̓�{Uv�CY�*��8�3>.y���[WuQ��#�Ղ��/^��4���J�!���Z+��A�����I���a/ߙ�����R�l�e���>Q�����6��,F���m�h$��6�,ݘ��ш}v�j>�."��$p?�.D����%���;��m���=��T�䁻V�܅���V����:�JƢ)�G�U����e�=~E�����a�#���U�'��>q�NF�na,@��1�D�?6����z¸N �Tc%�U���g�poB�����ϱYA��V֓����ay)b�+�����W}�>j�U�/ʿK��4�!jGG�1��?;܄�ɑg��>!���� /j�'�&�p�ч{�z_����՞Y�M|E�|�ɺ	����K���N���Jq��g�$��p-��{�����(#1��S"�"-��Ü�^����,O�&#�N���z����j�!-����`��e�����W��=*�������%��|�1����k�W�����Xv���ʪd~ނ�-���A��$G櫉�y��]�����W���0*1t7����S{|���'YI��&C���|�H��y�y9���=�OΊ�tG=�aQ1�r�޷	b���a �e�'�c\�����u	'��I�%�ѱ!��
ǡ�ŒT�쇈����ʇ�Y�x6B̧����C�� !����+nPq>�V��U��V�N��m�~]Y����l��¿-�����փq�H鬩�V*��wcsӮQ>��/���\�&.�KXᔬ�h��28��z9�G��L���(;��p�{6�}f���J�P�D�_��q��n��T��~��j��w���PFy=�N�e:�R/)_�ald/i�t��[RQ�{�3gS˓_{:0��f��wP
KΠ�櫙��������<�f�|�7�ntDD������|�"��Z��%a������#<�s�
�EG!�
�#����k����LP��α\�]�B����vr��t���U#�c�h%K��U�.�Wg� �Ҥnw��C`I�b�qَ�����'�w5w�C��	���։��C�a'e�dL�&P�#��/�Z�CӣU��5R�db'��;S�P0\W�a6�^�*l�$�Yl}�$8Y2Z%�t��PeFI)9�$�z��$��}��a7.�}�`'E���M̿��|E���>��.�h��C�������N�����D'��ܧ���鏾�_�9�j�g�h���}�6��;�n��Ƈ��"�u.��w|!Z3��{ ��@�N��9?~"X$D���Z��Z�߆�*��T�a���� ��#Q�>�8s�UH�l\����>�H�ɒ�%�d��ߥ� ������?{�����<7D�jW��רCv#:���طi���)2���_R�oP���=����mnC��Q5��[�p����w��slWvE���3�]mο^]�� $�!n�mg��c���e/��j�\�|��yD,�+v}a7�^�=̄�������� 2�+��y�ÂM@Bss��f���:�����D�]�L��?O���mMur�e1�N� ��q���\k���f�#�j�E��E���TR�Pi&��\a��!���]B�.z'� ���9q�B/{]q.�=N& ��å=�����������_7���r�A��"�I���5���V��a�ǻ�lǴʘ�S���^�*�ȅ3����CP��}�8�/a��07�{��_i���&b��D4>�˜Z ֡�+���k�!������ř����QN��A�@T��	��"(�|�g�ͩ���;/щ�dԯ-�o䖒��H	���]�,��l
G����R(����Nd�������lI��,�P���x b#��'AE�09d�w���>M�y��,z�2��pl�>����EM���V@ęrqъ�ʶ�p��!&�P/�X��$$Y~��y>�W+���=E�+��o�N�grw�/��m�`g������Or�o~=����I;�9��7�)m��7�*�@��ߞ2W&q��"�h�o+�ׂ*j��c;���}�9M��7�x�5���<��N{㵰3כiOr�{9�]��e*�W�|N���9��_:�uq�����.щ���BQ�g�\���̠M`j��_�a`/���V�)������������GI�Q���������6\_o��!��eۖAY���x�����w����TMPx~���)�z�p����Q���FU�o��+�W������5,�9�<x��Lu����WQ��
��(�=B�:�����CN���������C�8��M>LA���rNv�3����bL��$W�oqe��7�-�]p1gf#�u����'7�L>s��ô�S�OͿO�[Ԥ��E�̑'�m�P��A���j2�_�[�"">��J �z.��8������h'��'̯{��.\��[sfi������4EW�%���N�ׄ��j�����M��P�㿮���"*�d���
�i8rU�`@� &5l:A��w�H0wB�뾨q䥾C��4�}� ̣I���Nl��-duY��d���5�g��oX�qf��SP����mY�$�4���#b������Ag�Ҡ����l@w��$���`&��v�LKSor�h�0��5���|��y��'nd�4��Ύs?h:��\��
w��ސ5>�?�N3���&9,�$�w]�W�5Z�
�JQzl����!��D�����������r��@��K@@$�9G@��Ff�+C��(3��`7�wnF�M9��6Hp(����R.�<5c� =o�"����$��gr���F��vȭ�x<J������2"���9��j[Y����3aC��ܮ&�&�(+�@��}����Ǎ��s��]��j��q@��oo?}NYm���� o��5r[}�oO8�݄����s�p��u�u�g	�$hK?��:������g��H^p�s1������R�*�Ն�M��!\�k�Jt�JD���$�*��pX�b�"�T����pt�uc:�A���w[-��trA����L�Uu�T�������l��N����Q�3���"{l���̍�k#��E.8����$㇙�eX�j{���K@��8^��1�x=Æ�%p�b�s�e��X�ݏ��%�����b�Fd�g�G$q%I��+-ڼ�gh��ѝB����=��ۦ�v�����-�zG��$��`���-�j�.��"����.���&wzWG�J�W�NJe`v���'���
���B8^nA�_�>K,E���R�jedk���)"Ög�Z4���qr@N�B1y� H�����R)>�"p���i$�8�j���H��Pg��@���{jw:*_�y��?�����뛚~Lv�C3��ݿ|�$��l�����1!����Ow�O@���t�!B���sw���IKaS��*�I���L@�"�k����ۃ1s�u8|���O{Ro�~��Js��q�ϔ�],4ū1H�:�#�E�
H���%/��I[�����g�9�֋�?@�r���?͓���SN���!L��E��z�p�3��oj�J�d�D(j�j8m+t��Hv 
��WU�ŵ� #��(��|�Ue7m��@���]Y���)j���p�o����LPYs��7�_m)?��$(�b�?$�v���n���j�H��l�˱+r�X+S]9�*�z�`#����6��i�U|��C-�a����?��c�L�^��T4K�_��]�9�%���>(����������;w�N0�1@��}��孧��L�i:fd��A\Q.�-J>L' �po��נ�)��(X��ߥ"���:m�������Yy�Ye>K'xՓZK���KY���#��]q�VN��E� ��;|�Rm�ޛ�:IYٳ݉���̊o�P@`�d'k��廛����rP���*$��>|蚜O�c#��E�C<0^�_*i^�c��:[j�]��\bD'�"%Xp? .*�H���8*U��+��Rfb�MG�å0���Ax4[M �G�A����2�h��P�~��HO���.\E��{��d��	[�&����#%�<�A�J�z8wmf��X!K�m�K[�%�/P'�qq��$��mw�a�[��)^��hm� ߭�<Ӷ��]�D�2��Ǚ̆��k�=���>Q��c��zX2�t� �j{��xnW�E�^���#�i�Ù���g<*9�X�xzO�B���b:�Bk%��V�WM���/�S��Hak}C� ꯗ|��YT�
�X�&\�G�ǪU�'7*�m887��P�-��a�کl��1vDr*=�t���#,��;��IՍ�8�{p��}8{��K3T>�o�����v�9�F1�/�I�Rx�A�v%�A>O��7C ;�?2���)3r선��(�oᄸ���NhN���?������������~1�l���S�h�/(!�4�0Զ����%I����e���v���j��dr���.
��5�DlG�x��&d�]���	��jY��ː��\R���3@�*Y�m��nU�  ���//����;'�<1;jT�
}P�������T8ٸc|��(�P^5����&߯m���z��C�(�2�e�R�c_�՟�n�,8E����@]a���g��B��ۻ��&�7R�|<��(��,�U�����ͮf�G �o�UYp�^V�cC��u�'+�^LƏ��#�c.�)��Ĩ4��ϞE�E����w����������wl���c�m�y�~���yz��^7�0*��8�������1�&��#��,Q�̊?����G�B�߷��{�k������M��M	�'hd�V�4�^p�nY@@&��������Tb�R4Qzob����+�Ih4��M�����CV�	QP����Z��E��^����ȈX��a��������3�
ب�a���|+1�O+=}5Y�e�L��"м��=��w�H��j�����^��{֙R�'g�%�'���u�m�N�c$	T�k�O��¥���p[ᓡ+�N�_�==��c|h��o����^f���+(]��U���w�l1���`pL�������3T��75�2#� � +q����b7�5ڷ[�����oG~��A d�5��ǿ(6�����{����ޜ�$Ώ�؀=�p�3�Yc
t�w5?e�h�
�ܼ�~�6u��KQxo�4nwНh $q����Pڻ7Z���`r���-��t�S_[N�*�<q��s>Q�����J���t�[@����svi3P�#+���6s�7���7%��b^_7'�8D1D��Lp=���Z���l�+9b*���Ԍ�L�h�츭n�H��k�U�<�<.��C21�x䆡�G������(��^�3�Y�$5�Vؿ5n�sL�?=~�!�~6�eFJA��l��ȳ%b:����?�rM��d�S���l��؍��@P��m0!��L�C���]��%.Lbb���΀#CE�M�{�b��¥�y��w�.$��0�R�EJ�ώ��WH�i;��`u�k�y�BW�d�Cb����JZ����nR�~D&�Ǽ%2"�����/�"�j���X�*m=�A��q%��V����@`�(u�o�������7�O	$��^����������߲	��(��6uo�o
6��k����խU/�4��,������$mU���\�F�2�����Cl�pB�D�V��Z�⸉��	�|!(��7 ����S#�"8q�FNBH���+&D'�)�3���{G#hE���������@��6{�i������5S��7
| X�p�R��
fȐ�=g C
��[��o��_���`"�{�.1)8���TH�DRӆ�Fڱ#V�m Q�_�	����s_=�us��� #�zI�A(���;��G���jSvz��M�������ט�2�$s �P}�|$�Q?o~	A/�Ql3ⶍnь6�������+9�^$o	�Ⱥ���Ժ\�p��<�<��[0��)?^�X6�6� ��eO��KKtӿ��'1|����F����T��FX	'�!��b�;��`&���)p��χH��o���������3��j�a8��=w�n�ͥ���s���t�O[̢���U�INS�Ї2�q�����.+B�����le������w��_�~l��h�\]=wS���m�������ÖOt���S{|��,����!��>�Q���y�H�Qֈҷ8Ǽ��O9��������E3�.�̿�h�ِ����`��*gw��k1��`�9��̡(���<�I���X��E�aOiv�r���G�[7��]%x��8ڎ�ɼ/�yE����M*��\778z�ȗ&c�1_�/��������a+��ji`6�LJ&7弪Of��'�r-=�����ǂ�RλR��~�5�B��rŃ]���؊�0򗬲��qk�Q�6��� h�V\޴��W7z�S��S��.wL��s��L`-��Jp��_�f����>�Pf)��Y?s��}](f �a�\���i�}{���]?U.�Ud���%������/����s쎌��p��}�4�$߶�|ܽ����`�b��1
��q�ڎ�P��� #�ţu�>\b���a�A� �F��f�*m��e��^+���\����KK��'3�"�z������L `z�i��G�q%
��2����"V��T=i>�8f�}�<|L��6�\�9Bl$�n?]4d1���DIt�*:D���4����`?�ۘ���j�GD1mq�U)Tu�G{݊ӯd�"�,���؋
}W�����!�?!vsJ/��Sҥ��]�|�"��.��>X�����6A}A�a$R�KG����j��"���T,�8?#��mV�,�"�Ӎ�F(8�򶌬(�C�ۭ��d��AO��[�K�P�wNg|������"���O/���E���#�6��z�>�H��-O������y�@�}���M�	^�����.��Js�NT�<N( �
~�?��m�~��z-��g���Ñ�O�T]@�O���9*�����@�A�S�%��NzM�vx��FM������~	��%xք-ȞcЂc��c���}܁irp��/�=EJ�$�x��kCSh��N�u����F`� �p4\t��9�K 0�bkw1�3�ٱ�j�A���]�6 �6�K��߮p���>�� ��5�/�A}5C���ߐ"ơ������|�r�Ò���%�=Ħ=ƛ.�2�[�����������ℭW�l��[��m�Վ��}/{���^�������pԂ�/��vV-��?�  �5��+��n��L�s�x�>�A$��0��fM󪮎��v2���)I7�G?�ѹ�-BO$�Q{��p���j�-Q�d>dy��n[9�����E*���W��N��j<��j�~��Ͻ	��@%������Vu���H=����њ�$�Ze�Y`q���k��"m�N4o��K��T�C�����$��{���q#��� V=�b����FI�+L����+&�5�S�>X8>/���5�3�ӿ�ϯc�N�t����c�ׁ,�/X��X�x�k�ݢ��]�%К��e���@B 
�ys��"�e)ẍq�'HD�J��\Ѷ2�~^0Ȩ�V�$v�
Z���+�ea�يK���$�tH�(���+AI������[�`�6�^�,�,����C��ZU��*R��u�-��ͭ��?I�&���7qJ�����]��?U�_ E$�s����o~C�\��z�z]/�Nk'�L(�y*���4*�y-����ͯ����H�����ї@"�ZW~d�#�ê�.���"	)�S����<=2V)�+��ʌ���N@�:���w\��dn��#��c!R6��G��~��R@�No5-�}���C$: H�:�����V�5�b�����23���;]�~/i�Z���1�����*BⰞ�� �d���lg��Ĳ�'�Y��ų�o ���>FFA#Sy��ٙ�������q�o[I�mX�DOq\�ҺJ�<�6�0�p:��B�S!h*]A��A,��fɇ��1r�i�������jIT�uO,���*�=�p_�&(�#�mg�dX�.Ca��M�O����gv���5�<qO�=�g��V��Ir-�i�m�ê>�-��`��aM���ˮ�&���w���0N���Zҡ��s����2{���N���q<�Ob�׬|���ҫ�橳HvRs?GX
8x=�A�CK��c�G-Y��C�O<�H�*P!_�!�&���n^���Я:��HB ������ �H֚���W#�˻���:�����$K5�A��$Xh��ڠ���c_4"P�c�\,Kvۤ��醗�n��^�ﳚ��\{��	�K�7/�����;��'-u��u;���@W2e��!�����w�f�������Z0Y+a�u>��ZN���o��J[��7[�H��_��]��4��y�9�=�6����{�Ny�
����dY/	�� i/W����ä����q�R�Z
>a���[�<��J)��RTkݯ���e �ø�r�v�O.ms��/p�L�yO��h�|SZ:�!�0d�f�}޻��L����f�To���ݲ�x/o��|�
���<��˭�̙�jq��L�=B>!(	��gwn��`p�p2�k��}�I��n�{�I��4���sS�`�����������a<Nf�L~y銩
yoy����0�"o��&#_�`{����	��&H,�L���j�������S"K�=�cx{1�@�r�e����JX'��q���^7��T���k|�J��t����6zo�s��Um>~:���3�'f$�@��H�e�ڥ�:�L��Q��/��i�����OO�r١�ʑ��|�����˂�$�j���z���k�x�s�/ݮ����Q�����ؚ�F�[�R(-%��A�u���{�X���P*��ƖWw��Pďa	�@W��R����^9W� "r�`Y.�>�x����߳7��-��4T��e�p4V�����c.@bq怳R�X���F/-[���)�- �."T)�>t~���j6�q�]=����S�:�M/���Λ����`�2���&T�gw1���u5r��
r�f�ز�jx���xx\RdO^]��|0�1�;�-��'8��o�#�E�����h�.L���* �F���ѱ4�c�B�b��w�	��ߩ ����G�QL��.��h��u���T���L���0�N[l�՘6�R�+�>�x���A@�D�.&dw���T�rN4����@�tߠ��eN�F��~���R�"�Pq	h�}v��g_����d�~�e�\� ��.B�5$F�|'F���ϫ�!ɒJQ�1M(h-����f��^2����.Y��NO��տ-�M�U�(�
`G���r�B���o�f�T ���j��gT+*��"�MM� ����k������q;�Z������H����t�PK�,���J��+�co�P3��5����M���^�\��.p*�m27�0���&��ً�GG����a">^�2R�W�Z�>v�6j��������_�l:鸉�n��@ 'O�7�R��!j���8_�l���t�4،|�#�`����5���5�0�x��}�/�N0�O���_Ȱ�^�Kqx6�t"G��q.;��JB]r�<L���w����6�g���`B����M(�
;"cy,���Ǐ#'�������iI8�z�x!N(��O�v����#�`�p��֗�o��^���ؠP�~�ς�Z�F����;�4O�2Ty�v��K�����-���Q,�Ͼ\#����;�ty���7"�|F�x	���^��74Z���^��&Mx�H}�WA5�P	f�L�=p��B�9C������ꪸ��
w`Г�Hc����U!�$�Qz�#Í	�Rg��~^E�o�Pt��K:r��-��^7�b�y!g��A*sG���R_j�E��Eѻ"
��r��0�8L:]�X�L
���3��D���R`�p��ף���W]��>;MHG"e�p4}��0���z�i�V�`�iڑ�Gd�6.�ދ��B-���"�J>h�����<���e��b� )��~�1uɥͭ]���s��
,e�h_��Vj� ����	��d5������}�<��NT��es��Z��k�58����.G"<��%���?��]����x��~�72�"��o���`{�7���� �
j�������-�A)��Srz��}>�����p?SVټ��6ç�����-�o�[�>ő,�q.��à�/Tس�X�3R��!Ζ�@i����Ŗ<ߎ���X�u��sdl�u^�p'0�X����cL�Xt��mO"�`�]&�x������MJ�d���ep>��TֿG��,��g���]��@-r
�e:���Q�`�L����H��.A�������1O٤�M�n�
8��Y�,9x��� s
���
�,���8�h : 15�8�Ts��,bn���ǟ��H�b���p� �3���ĸ�����q��K��`�U}����j��Zf�̎=�Rh�j;`Ä�P[�o�1-J���9V�����������t�����H�M����<�6N"�\��_0a���:cSo���� �3�r4|��\�(��q(�Q?$�b�6�;�,Lv�da5S&ڝ��v�)6S
�8�M�z ����5b8��nm$�ʾ_�6�J��aE$� �L&X�vB(��c �8ٔ����$�=������k���Ԓ弻:6�i�*�Y�jE���i1Rd�f]!Qd
��-D�l��`���ρ�:>�
wI��˄��{Y7S��S��-(=�;�_y�Fp����2,�e������]�ww��@����Cpw���Π�9��{����յj�Tu���|ָ���Prצ^��Z:p��c� ��C��ߘ��z�,����C�A���>��I������n�y�Z�LKEFKI�-�.����Mџ��(�H�����ǫ7�GJ�{� *�����wq�����+���=�'���ԓdH0�
��Mӻ���m�t	���R�k����
���I�E�xr)��2���C '��R��|�	��u���P}!�E�#e����FQ�),jB_i�7���-����R[�lS�\�(��D����~�;�>dk~9���s~�a7a��[��3���l�bŗHSd
�ִ���F�SD.*<:@�|x����b��`Z�I%r�� �SY}����.�U}L��y��V����j,��^�
���J���	pc��^#�M���7c��`�ɺ��OL���8Z/�ѷ���.��ݱ���Cn�B�m��l��J.Ҹ��B��'���� _c��O?��	>��Q�-�+�����(6,��*EH��߰���w_-;eo��O���??�л�i?���XA|���#͝��bEL"<�XH�i������Y�0ҡ{�ɦ^)Y����f�>��5 �=��XinN#�!�,���.�
��)�N�_��v3�!�"�$T�v����@�-j|5B6�IEA}�����ف�������j��'Lh(C����$����FY�⥆�߷+X$��ӗ&�"��[�r敻�3��B�~�4��/���C8:W.G݆ސ�r_��xg���|GY>�i�8r�)#��A����=d�[U���39~��Ԯ�w��W���0[���.����H��*�u+�-�zZ�z~�
G�[�I�Q��8��5h���ӻR
ʲ��{��rg�bL�5O�������+)���Z+i}�s�5w+�p��_�C�}���2
�n��DɕQ��L�.y �_�����+yv�^��jl�~-E��& ]�q��=�\7(;�j���Lec��!�EL���-ȍH� ����H�&�ϊF��_vs{--0IS�?�w����:�+?�k5�&�8�|�O�o�Xh{v�`5��p*0�uf6��f9_�;�\Z�3����:�������9��t���\�t�zn�R�\L��h��l/3Ϭ|�&�� =���9��l�]�`�(�P�w�F�KG��dL�Ҽ�Yz2rK�����)������ �Wz�cC���/21�y�����T��<��kG�6�ʈ����������!�d�3ٌ��X)�B�Qf�>Cm��1C)��}�h=(Zm����- ���&Bu�Ǌ�)�ϛ���x�xW->��3��T/��z�}?Jdh�cEԮ���@ߚ	�Uw�iӺn�\}!�db�����xRR�jJ�I8MA # `�m/���7*���V�Z�F��&I[ӕ��;郗
�E���8����P�
ь�!X�u6��Z���C)(�	|�o�漌C�	^JQ�C�>- �񀏄�8f,[��}�E!B�Bd�FD�*�b��} �H߃"~�-B��\��7�o�R\.�-bξ��󃍛������;���\}p��w;o;��A�0�2�U�UM�D�����i�҄�>f����������r��n!��߰R��=��t6�������8y1�@����h7[qJ6��z$�<���DBGم�.�>O�˲kw���+UWkyk[�鲎␃1jEДΟ��%�"����q��0�2	*A�5ܹjP�0�F�Vi�b���󎵾�[-uw�^�8:�_y������0(����,��	[�Ȝ����)�ehe�i4�z%��x(w�xym�Y����t"�Zq'�~�^���g�� ��B���,v��D�W�h�,�ǈ�U���W�7���$f���Kۑ3�k��J����x�x�������^b0U�c�	ɇ�ⷷӨ�d�E�=�l�L��w�, ���G�0$�4zn���{�4�)��.}4��z�ۗ��kw�p��j�)������l� ��*���յ��:L����Q���пRbҠ/:��\+PE>��d�VԂ;Y��ꁋ�����ϙ/�i��brk��
�]�C}�y�5U�Vc�k�Yxh(��Lv�*��߯�s��V ]�� �� K�m��#t���Fg��b�=���\e�S�n�'�誉�v�4t�n��&N�IO�����B�ЁoJk�U�5><�h�É~�+����njK�lQ���ξr���7p
��OPO���Nٞ7i��<�����8O���&D��tS�v���\-"��48<ˁ"�&H��L7�1��ߤ�|�����RlP������*�A�C��F|��}����#X�h0 �j��|wcI�sF����UG�Mg'���x��j�a�חh8C�/@Az�Qcv����JZb��t��Ϩ�+�{܀Q�X�C� =慤Eb��{v�g_e�jĔg{S�T���^�%��>JCV�Z�(�{�Q�Q��?��9�S�t>��T����1a��m�v���Sms���4�����9}K��9�Ё�X��fw�ZX[�y q_�-TЭ�h����ğ{��ױ�^�b���a��u�t� ��!�.�}��j��t�]�3�"�~9*�@�o1�X��S:�k��t���s�@��e�H��8�/���a��Dk�2���['/�^ӊQ���b�AV.�:3ı��;
�=���Q�*�9�����UV�^ج}�0�#����q�k��:�?n�_y�{���-�δ[iC����	�Z.(wd��m�H���E ������k��C��ӫ�'�[2E���U=.�M.s�Z"�{�@"�)��΃���7�8wbP��#�M{_� �)�o�v��x��؜��E�	݋�SFo�x���<h'���:����)M�9�J�2��4���b�2I�mQ�F�Z욨��"w脸d��۲���<���y z���R	�����gu���-���0��g�;���FBfj�ո��������3�X��R"d�m=e7�t4RE�[���?2铵���?��E�T���_C�U�#�|V�~��'G�2b|��ҶAN$*J�(m���R���-�����	�'AG���+g�^�P�	���� j-����~�o�>�*Pr���o�e�"`d��yF�m�x7�z���u�HX�)c��Z~������aO|�$$3�
��O��͙��K,��V���>r� �@�1cc�����u�i�l�\�ڞ!�UY<�K ��&�roj�X]{9*�
Ð�n��3霕2������EQ�|@ 3W �;�2��>�\�����|�}<mD�0���1�'t��� Z��t-f	�ڏ=��v2s�ŲX$���_��22I�;�j!���b�	\�"�5�|��!����ʗm	�w8� ʍ`6W�4�?�n�棶���?e�+Z���;��)��A�t|�I"MD�#���M�-\���?_E��9p��@���<GB����}�͠��Tw��o�['vW*q�w䞧0Q�	6ẄIiL�vv���>w��%\� �P�R\��D�����q�B��R�[��}#��߉�~�����������M�k�L������~R5�B�-��
ϥ~/:TVM�i�8�r�;FaԀ���]����IFJT9�)�W�O�o�4X@�-1�Ly_d9�+��2L7YV�U�K�8Ӎ��������C�����SX:U$Ou^=�k��%hg0l���F���-{#W����@NOTLg~LT�>�$���J4��������ZȚ��'�V� ����!�<�f&c[o��7b�2K��ˉ|� ����jH
� <ޠ0�F#M��:�pV���ܐ`Ϯ�� A	%}e��u%�l���+����;M_R��D	���KjA��I�4����߫	�ž�2�K�#+�_��}�mE���H�̸X&b���ܗGi2�K���$��<Ī��3�i��Џ�JK�S�����U�%d����X0,���x3�"P#<	�15U`H��7{Y������zn����J����!y��b���(�~��b�Э�}�\*��t�������[iLM$�M^��I1��� ��6/�Q�1�ÃN����(�fo���k�Զ�)]"h��w��_�u��nR���3��Eti����f(��Dy�ŪZ ����k����l�q�+�s��������褦�U8��:9�x��H$w�xexc���GX�k�����̙��V�lX���E��%/Xp
mm���=���[�o�>H)�b�Lָ�8�Ų����p~?-�RF���?6���Y���)���nP,��B�ʇ���ngj^�</�]
ʺ�aa
�k�@�w��2/��7W�M�����L�:آ���p�ʆϛ$�}[	*Gi�t�+��YE9���O�>��!"�q��[����e�ڽǂ!��D��K`�������0���ހ��O��X�Q�F�L���$�Seb��9�p �CP�w���ꌜ������v7s�O��au�kꍻ<��6RN��%2o�nnd��"���%+s)X�S�u��F7�j%�$��W{�W��T��:�`�5p\~not����h� �Z�I=�:u�[�8W�<]�]�cS0L-�T�B�uP�mu�u/w�o�뀮M��s�P����[�F�x��~;jMG?����-��{��-'A8��j�Q�>)w����W#JW��\̀PN�O�Y��$�쌈�=,���Q��}R�FCk����/�@,Xus��s'�%7��D�?;6�C��%	4	�I�\��`S�H�*M�@Nb��x�U�_�9J�IDYy���uO��駽�[���G:��rE�����WW�gh&�C!Y��������V�{�M�"���$^Z�+���mM_P�)��:Rik_H[>����r�*�?��6Ń�R!dzq���{�"�q���S{{9�~lII�<����_x��t-�yO^Nb4[\��sc��B�.6�~����W����E��M��o�=ۦ�p�3n�Ǭoo�$B/��pi�Vy�ï5�d��*�O�}+�rx�@i�-�O�T٫�FJ줪����_L��
����p��N0����=��PR ��@"f�vü����9�>t�5�pvz�g��Z���b�l����^��E@5[I�_�MP��=�CW�?�D	_y�G���]�a�?W���O�A�}�N<��^K��@q}yƣC����L�*�b��$[R���y=;SPN��ay(���P�[M^:�=�\�)����@�w��B�<

c��]  n�"a��y��{b�_Պ�J��F�ͪԒoE���:zk�x�6{�=�{a��j�����%���<�^�O�)(q��.���O R��3<H� y���nM���m��]�~iŅh/9�+I-,�:�a���f��B�"�3���$��k�,���,��9���=��]�?:����DGKkm�j�!`%�B��H�p�V��IjۭjS�L�ށ6����(���~�����ڕ��h�n���B�e���oG9�d: 4�=_�����d�"�AaRm�=��%�M�0����Ҋ�6\�
�7���d�^�7��Ċ�Ȗ�� ~ � |�P��\�.�"n`Y���Y<�x2¶.����+�|�ɴ��}�e���ѱ���LMp��k2J� `:qZ"s��E�X��M.a-y����x�\�7=me�.���ǖ~Iwn���S��˿��*�*�=*�G�T5�|sS��'sNLr��}��ZC�bλA�S�
�G4 ����tg�� N-{ޞb��Dd�j^�
��rHl|�jӦ�/�M��>AF���lEm�-9:�Bg��`����Ţ<��H>��$<��։�#�p��m��&��Z��<�w5A���R=қw�iyn�2��5DC��E��
�E&������A�%����7 ���FB�[�|�j�����w�
�3�{EF/������j+�� ����`�AL�	kEEȵG���ʔ��ۨ�k�*-�h�j�Az3V��rr�4�r�)%lp.'�|�Q�?֌���e�6�brmI���]�<�%�A��7;�rݔY,��x��5�ٽe|���%ް�궍p�Br�n��0}�'}��(ϵ�"M��y���3�i��Zm{y<��ğ��/g��뺓��y���H�]�.�d�e��r�&�fL9�,zxQS���onL)�.R�q��>m�c״������1@��U����M��M��G�.�lp|�P�����ك�h�f��E�� �xY���������G�f�����E6ڒ��poz�3ͫd��`));��,z��!/X� :׾����}%��b)E�
���{7v~�n����9�}�#To����S��n�����2����o���+a�+�P�/z�'6��Rt�x��%�C&b�og�u�r�@�އ� �%'듞AN�f;5VE�5_#z�;�9��6����O�B������Ww���RE���l����EɈ�Bc+I�'������r?�}Ӎi����дǈ?%aj��M��>n�&��<f�Ǩ��G2ÊDj�	�D���:ɪ�ث�%y3����Z@�͛k���#Pt���x�=����<%I�诋llN>='6〦D1Ѿ�������^)�Cw��_�e�5�Z���V����{��S5��Ϡ��ʝ�2�����O�]'�������^2�������Ca��ᨸlf�*��X�A���=�����;�P�T��q����g������V��T�/eM���W!���BXϥ����x�4,9ۄŷ����dA$��id9x�q�	)`������]�jG>�'*�]�t�K)��KO'VuWvUەv�(=�����_����-R%N��X���"��ٗ44!G��3U��S�FS;ʧ2��աIឬS�9��o+��jf&z�i�lo(��X�$�7�@}���^�p�'���c�AxIgArJvHXϵ���Շ��u��0}�]s���%'el����a.���T_�<w�~��J��[�;j����-����7�"b�u�VZ���+*��-G����x�U���+�.�=����~���;���v��@�W^u0�(�@Ď�kL�LG��s��:��LIB
�tu��W�j�8UQF�;o���c̮�M��sd��<i�H�`2�6+����Ӥ]A��i�X㟹퓣_�I�����6�v�~k�^,�����T��8�9��cd娌�%�d��zDU,�x���O����#��Bc�	�q��~�.��,���_?}�RH�/�Ϥ K��:;��)c�]�p����@OY�5{�t����;�2�!�����߀n�W94��-�|����y��-�siHEm�,���'�*x����HKH�^Wjeq ��hV3f۳l���r���-,]ŕS*�"u_�D�!��üx �h��*���٩��Ҵq)���4�ЭY�"ȝ�� �W���D��[���`H{�0��&���(�'���O�iɭ"<��-�K���%�����=[W�!^bS����!�y�c(t\�D��Ǜ����o�e��dJ�ru���/�9A��C'�*��<���8�\ٛ�� I�.;}���?��N8�J��
.�]����J���-s�/`%��+:�^[B,�_h�+�ލ:?m�}!��0���Ig��~˟�����-�.�S~o��,`O�O�˾�-��h���h�S����V���&M���SsZ���)�A�|3<.�sb�R�S��׈q��ӂq���5%5�&KnqB�(${�A�6�K�]TQ>�������_=���4#�r��5u�@���r85Bg'�(`�C�D�v�ܖ�6+X������|���=JIns��Y���DV$�vr���	/��Z?F�h�da���G��c��eS���i�da昅/E��KnU��3�M��>���I�H�{W����
���(g�B�cp�df�0kd���a�����=e?�D�^uz��I7��{����h@��gٳR4��+�������2��S�9 ��tzK}��>�0T���Rz&�f;����o$�C1A���ֳ��H8�<w;��^<e����v��H��A����x/+m6K
:=�wq��DNԄo(
��e��&���-��L���Gp���2���u��1T1&�Xm�g����_��|�{i'ȓ�2.�D��x2a�l�?����}XZ��#��G����v�aZ��6�ؾ��J�)���9�{m��Z��i�����A�ø�]^~���)�Wz�cvj���s���垱h��r�H��O��~��� .�@D�(���z��v���ɠ�Hijx����։��w0cf[�~�Lw	���`a��J�(�M�e#�ɀ��S�G�b3H3@����3�zLI�~���/����
-kj�^p|mvd�gIO���\&��Ѵ����T�W�l��,b<G��g��F��0�0���<'�N��8P�{��sm{���ٱG`5ԭ1l��g�&%����U�^�-uLII�,���J�����4����o��͋"�G�l��5p�C1���>�����"Tu�Z?e�,7��1�0V�/T5�VR
�FEa��~�������-Ծ]+.ꓐP'f��N�Dw��������!,��-����ex�Q&)-?F��O�* ��P]?c{��j��l� <m7Gt#�L��G����c�؟�	$hH�H!ڗ����w��69�W�Ȣ0���_H&�ަ���"���b�H��L�+�'빻���gJ��8^�G^;t�j����{	J;��7���� Ot*n,� �֖үH�@޶�M�@@4�éX�.Xܾ�?�N��l+s���^��	d>8���6��?��HR�sB-j�Y�V�u�B����D��%��,��T��*����X�x������r�/b���^��S�Q���4�?PK   (_�X�����"  �"  /   images/83968c91-e49e-422b-be2f-46fb404d4a04.png�"݉PNG

   IHDR   d   7   ���   	pHYs  P�  P���Dm   tEXtSoftware www.inkscape.org��<  "pIDATx���y��U��w�{kJ���2UBI !�DA"�Jd��->�x*v�zK]�G���(�����2=��L �		�TU�JU���y�o��w�͗�M���֩���θ��9_L��+5�W��5G4�(����e֬Y���&���RZZj�g̘a����e���2g��:u�����Hy�AY�`�L�8�ʎ;&��s�9GƎ+�x\>l�K�,���+������r��Jn^�h����K�.���l-���2�����;O23�dpp�����om��ӵlP���csg�h4j�w�ޭm2m.�HTzz��^nn�,\�P�G�����7N�ϟo}���[�)S�HQQ�����ظ�=��q�����_i�s�|[��ͺJ�� �	F�1a�1c�Xx�XXɬ�l�S�Z=RQ��Sh�Y0i޼y2~�x�q�+�a,�z�@���@�!MK"��ŋ+���l(�����ٸCq��r��u>�A�H�,[���g�V/-.˗/���?''����͑��?_222$;{��5//W.����-�YY�V�H��u��6��q���0�4wh^�ȟ�|S,� 2k�]��!�h��Ha�X���%S
��92a���˼	ݒ�5$�+�����d��.�Ȯ#AY��-��)]})�ɲ2ڮ��!�m19X�i���ʧ���PC�m�P�e)%ʥ�ڥ�:Kꆲ�3 �guȎC��8r��䳋:ek�rNN�jж�������dDe�y�,�
D�d��9]��4G;V�� �O���7��w�ebn�O��AQ6��Wf��-�y�_(=��_5�i^��7���� �n��͚�I<7�-��5/	) ��7*������D�o0�T��֮���2�5uƴ^@�^������ֵ���j���?bm�,�IMkz�����ֲ�����BY��,�+�g�2AE�����o "5:n��As�m�%J�2��О.i^���K�!�5wiި�� d��r�[���G����$��:�|i�[�Uy^.ӦM��h����`��;Xnb��=���w���#2{�,9�:���z����c2w�\�l�1���*55��6�8ioo���F����ri--&����V˴^CC��1�YiM�Dӆ���Z9k@�2SJj2$�KU�QC�4Յ�E�ޑ#�U�d��)S���E����$Bt�$�W�ieD��r�.S��7��G#c��[��1�d����	F8�yn,�f�k���>��!uuu���ۍu#
��"E�¦(M�켌z�nkkS�5����ߔ�d�e�_6���@�2�eMM���!�������̥������˨G�C�����{ƟX]ce�G?<#��GOOOr<tW���ѣ&j}��-�&� #�7J�%�5Y����VF�CHk֬�ɓ'KGG����UV�Ze� Q ```@e|�TWW�$���.��@HXO^x�!�	�J�-2�����I�&Y�|�)}�0.ϔ1(�� ���\������A" ���!��7s����&�qS�  �{�����ߖ�+W�a\<�����e�]fk���\7j~D����I�OwK`�"��k�O	̍*!> �۹s�Mj0,�Hʜ
��ar��Ƃ $�c2��ȑ#f��t��2�ji�����Y�����7�'��(q�5sչ���ː��/c�y��qP���q*��Oo��:���3S1�ܦM�nEEE���jY�b����R�|�4�^s��F��!P�W�u:���L��
۷o��3eήd8��x�y��7�>�#C5P�@��:~�������p�|�W�Y+�Xc ,F���Ha�!��ӧ�5��HΘ,��Ҏ�"J }:^�X{z��6����+=�u�$ѥ����1ي �'��I��ի�c�b��Ա�y��Ek�_�D����3f���
���?6?�#e�	��C�i�o���}��GM����ʰ>J���/���۸��;�AE�����7��"9����p�O�[�t�\��+�y�����wݩH��}�{�$�.bq ���A~�ؘ������Ųt�4y�߶�u�_&ͪI�n���޸B^���5C}����?m��CG��l_������4�c�{���d���!�Z>K��@��v����Ȗm�r�Wj��2sz��9Y���۴ϕ�g����������{[+����Lfj�Jԉ���?6j$�%�s�=&b ����M,̜9S~������G��&s��G�'D��wݭm��&�QJ�ʯ�_v��u"5�Tt��%tx�������,�}�.,6N����Xd��=*��&���ϕ���R~4OV_|��4E��[6WJFd��OwTT���k��õJ�铤���RV���Jsg@�\8K�VFd����{��4��sR��}Α���[���5Wɡ}��}KYe��_����,+�!b�u��OJ�=v�%��ۏ�裏Ј�;�cJ�ӟ��a��_V�8 /���YF���Ɔz�U t�	n�K�n8�O�K��3S��ʄ��f���~e����}�����O��.��⠽�û����uލ�=���$��=	`"*r�z �y!=H�"��$�cP�"=���Fl��,Dy"���S�����-]�0�"LsLe�Ͽ�zx���G���:a���z	�7|\��immI*g�h�o��v.&�/��GB� �caڟ��C�yb{����3k�-��w�}��)���@�m�f��e �o|�V��q@O���$bS�'��S�k<��To�����C��M
�瞓/}�Kf����@☄^�nD�y���Q=��w1�aEbQ�j3��wl#���N3Y�.���@F����{fـ0��[o���r�k&e�@��{v�R|4)6|�,��yHߵh6��ON���|��&"`�c���φ����7�h����ȸ�~�/��3�! ��'HÄf.�f>�"R"C�B�;v���b���$wn�'i��L楗^2�v�ڵ��� �I���!��#����Sp�#�����r��9�%��O�ؒb�b�*����`����ȑ�!㤫���l~2�""��  Y����(u@\򤓉6'�A_n��;iw*.9U�.�z�	�|�<O�x�(y�q�7ʖ-[N@��Z[Z�M4A���:��T),��|2�7����(0��f������;ԏQ��tu�����7������%Ͼ�S-���7s[�bE@ڎ��!I�S���snIe�p�W�g֍�{6\�8�H��b�' ������N	+'�`ee�Y6tx:�6�������֜�C�u�2$��Y2�S���x������Y1ɻl����͔%�L5����������N����l�}(���l�aY҇��F�wR2�S)1!懄>��C�h��;s$��ݻ��S�?l���g�Z�H}�|[,Y�Rٻ���d�6�ʴ�C*͎��<5i�U��7���y�ޛ�`�&�2��D���@�H��	�aU(n�!�0Q�D\��[��l����w�+W^y���]w�e�qx'��P�٦��xA����ʖw�J���7�"l�|���Y5�ӓ�R�ψʄA����C�y������1\<:W����b�t��[�\����l��C�J���|g<�C-�9�ǽ��+���j�!N"�sVu���Ǩ���=�|O(��UY{�W_s��^u�������;,+�Н��e�ª�ќ3g�\�z�4V&�Iy��/��֓Ň#���y����!��I������APD��r��>����5����o���f`�Hxd�.����c�=&�<�ƫ���@�QW�R�u�� ������G�(�w��Gy��-���o}��ҧ�xB���ԔdKK�E @<2��k�Qjk�l�K�_�{A��X�Es�X�����"X���J��,J�p�ъF�<��~��%A��g,���k��`g#��<g͞=���m.? Jc�@�G-	0ʭ���$�p�"s��0�_� ��hl��Y3gK_o��< ��כܣ�@��nQ�l�Al F���l�ٛ�Қ:�d�x��a�A 2�|
�1X�w$?$�:�ebD�;� -�d�B/�����
"*�S:q�m O�`�'f{�j�q� ����=��s<^��,++I�8�)/�/���V&��cǪl;��K/M�E����6�S4�I&7� /K��l��Om����b�X4 eN��7z�Յ��b��aB��d��1@8�t:��Aux��
s
	d���|�:7���e�$�D����d�V�ѣUI3��VW�Z蜄N*Tj�8X����d��ܴ^������7����[o��a^�r�/_&6�ju�;������3�N�p�U��&�5B0�SI0`�.N|˙� �}�T��$�J����+s&���N�?��(2�Y��e�I"�W���_�w� ۷o�쉾���O����ig�%N��|��f�r���O`7�A[8F֬�cGsR%��C�$c8��C��������Ɔ���$���Mo��"���p���ş��v�|�o8�	����roy�Ώ�U�O�+�/��[p��c�:���t�=�q�ֹ ۴i֗�+_c�u��t=�&��0)��t/��(��S?]����yx���.� r��jY�l������-e�?���vp|���R�|�9���9���w���,��}���[! ?�;�ԁ\)�� yg�|�s��=���w�A�4�L֭��&WVv�8��1*�6�i�k�~J{�{gg�^�[�y��4I���7������:��ks��3��;��9pg�q�<:aTd+¹�x��K��͛7'�x4ł�,���<��}�D��L�l��T��$'�f�d�o�vB9�[�Α���H�����2�x�)�;���'p�w(���c�9�Q"��J=t�h�*F�4�/�d(���r8��d`s?��1 � y��ǒTw�Й&��c�G���N�>������ma���+�P��$Qq�vJ(yp1,
InR;�����c�vGd�Xsd�i�h82h�E� <�n�р=j
`38,Ɯ�����?�`�<|�� ')';C.��Hj��)ڧ�bF���F���a��uE�}���i���T퉠�E2<����pVcS�mK,�ܕ�P����'�|2����;aSz�D�I�&���9Ë&!68���IZ�z�W���k�R���&;'�޸�''�ᦨǲ\�x�NH�|ox�c~ZнW�7my�@��k֬U6�ׅ֞�)�/�~?�����s7�f�IvAzkk�9��p�4_=�u�]$-]�ޛN�ׇa��u1w�+e��.p�CF���ew36j;6H�_����P^8��s(�M*"�L������{v�A�+ s�z���D
[r�v4	J\�r��;�q,Z�0����+7�؉�R�� W8��)�Bq��8��<��.�8^x�tɈ7'KV�?_j�e4����z�'��)w��_������?��IC�"��X'NYpD�#6n��qԁ�	@�N9���Q���S��h#	MS�(5N%uu�I�F?9���5�u�p�D�� ��!� )~P���x�D��� [�.�-o�,8/6
��@wR�?��S�?�)ɞᐃ�w
;��q��h����'���������@� ��������㔢�%��+/�T� 0,�����\;�0<���{2��c1�`��	XZ���hYă��ڜ�FY�>V�,o���'M�'l�~���7���w�5'	������<��AO�cN��ku��w�<qB}��7��htPuG����U)zlR�q�=56wʿ?�S.��̓j9!��9έ�(�a^�Dc Ġ���)���n4J=pF�k�)���ݵk�\q�F�t�����5�\m�.Qx[�l=#�)�Pf͞m~D{{�����x��\���QnzY�1�LN��\�i�X[z��!���ALn�;���� ��p
F'5c ����j�(����Kd����M"䡇2d`��s��eQǘ$�w��i�=��W��&�1
��%8 44DT�u��2��	@���l�u��C�w��a1��@41�v9q��n�l$���W���XuHը8b��2�@�'�Һu��.;rq�%r��!���{F���2}/:g��ٽK�[�%��(CL�TU�*��Y�������"��&I{��ɣ�Wn�Z�C�xh�nG����{�X[��X����ok�-�h_]�6��i1����O�S����p�5:{��g��?��-�@)sWJ:��/���"�1���{���;� i��-v�=��E�{����?�)�o��¡?�@�D��?����K�ͪ�I�wt���XnW1�.1��a�bU1�_��I����nR�q�!fӦM����&ĭXڀ��F�|o��G�\�`!�`�V+{�|b'T�9D��ܹ˨������O�: ]$����Q��7s�-��C� <��g����X��Sb�.��q���+A7����o$�d��#1���o��V�����0�pi�3�''���	����GW	�p�ȯ�s<�& jZ�����͕g�:��񹤧�F�?%B��v,@�'�}h(�Is_�|D�}���ZX��@"J�;(??��=�#����T�`�|��7n�h��������0�&��S�T�2���|��=	 �D�'��]P�AL�Y�s`<8D�!�p�� �."}BC�����{��6��k���g��!?�я��1 ��<|���;����H8�{��N��wؠ ����C�	���loo_�T��t�b@�7ސ@x�!��U�M�v�r PW�(����%�䉿| �a�46u��ͫ�6|"3�Ȣ�)��3[e��n�:<$�^�(��fI��,������_]-7�ܜ-�-xz�����-�o�{���������3�d��VG�to����er��.�Y�Չ�hė���n��6�Ǯ|�~��X�'�0�GM�{':�`g�> �/��5�T����-�
k$ l���u���޶mۓN�By��]��;�j��˃m��m��?����v�0a����N�R���Aff�|�����I�1�m����6$/m|��|����[�hlD�}`����+)���7�R��ȯެ\�f�������]}I1�KB-���C�9�湚�Y�pe��w���I� �.��rS��^{�Ev����N��'f�肛� Āg�t�����17n�`�n��H�\gN��R�!�T�}��_���&ikm��7�r��|RbD�q7�Ζ- CgaX@$lJ���{���믿a��H�K,S7|85ÁA��f ��LD�2��/7
�W�O2q}�w�S��$���<ŷ��~I�fͅ#a.  ��t��������"���I���Y ���=�nx�׌��N �{LZ���C���m|%"8>4(�� �4��-��Q��}��Z��BԀgNUr��q;:��q%��z@
Ҁ�p�K��bg{��PX/D����`�:͉mO�7�e��!�X���apFA<���i�����|�t�Ꙥ�$��&
�6l�`�P���2Bh��X< g�hD%��m0�$��@,�F�S��v?��~B�2 J=?�ȸ����pm���[%�M�Dz&�OK�i�)�!�Q� M��� 0�{Vv�����^�ó�se�v�.#3؛��갽DA4=���������fZ��tE���s����mjb$Q���`���)ត_���Civ�`p��ʘ�#,ħ���Iܔ�b�'M�K;��_����7]���\�!-�
M�ć�-ґ�"P*E��@r�R͗i~-T�u�	!�˦Ș��-c2��`}��� ���.��L+��]j*��R?d���E�T$�`N�1߄�y:����w��<3/N��V������A9gZ�mJ�±�"��i]Rѐ)�pf���Z<�[��f�$E�}K�xj���4D����H�J��dQ��>)��+%U�F ��̊�ɬ��R�e
e9�2�`@ʪ3�:��e�ȸ�9P�mđ@�?h��|#�z���B�@�����%�e��2�d�G�C��=h�
�b���w�xW�e�ǝ-��3h���dN4��Bz�^c����ײ�.��� ^`�O�뗺6��z�(`R��}u��?��`Pv�N���}q�?)�_��)���nv4��U�%����hB��/�ٸ%��\f,.�$^���o������˅�g5�)�� ��H�{;��[%�#���+�C|Hٴ1���Xd��c�x_m �"i�Z�d��Tei��F+�q$7�>-k��my|bQz���ݨ���|s���Ղ�z��/��ޮd�|���̞�;]�\�(+0�tuv$O��QVh�X�x��_�h�-��.I����Ҏ�F����2�^��ʽ�3[�;��Nb�* ʫ[���%���9�DZ�Ȩ��D>�?��M3����/g����PrX;��B^��4r�= KBibY��~V�&|���o"��!\�s�X,�CY�.�@�a�����n�����8��Q�E�B&��_%�9���O-R�a����e ��y��2��_q�Oq� d@����������    IEND�B`�PK   '_�X��iP  K  /   images/8489a8f8-4880-44ba-919e-53c698ce78bf.pngK��PNG

   IHDR   d   -   X���   	pHYs  0�  0�
�D   tEXtSoftware www.inkscape.org��<  �IDATx��\il\���6���vlǎ�8���',!��&*��@�JCKQ��O[Z�U%ğ��P���DE�P�hÒ&B��4�N�I��3�Y޻=羱�f�č3�`�|�yw��;�{o��?�O G�鉿��T
�,F��I��PY�Àl�r�|*G�T G٠f*+���`�0 T�T�S� G٢a���1ѐZؚ�R$P��"�P�UL�ꨄ�Tq���2K�S5xB�Pc�1��������d&�6
�QTw�3�	��,�dDE1��(b1W�:S����>��ē׉7�T�/4��cě�1�/�|�P,s��I�&����tł���;_�2�G�h��
�x�I�A�-�-��ϖf)f�fŊߐ����.��
	�'�<!�<�'H�Du�����~���j��f}�k+z����U`w�
��^��;K��F�ŝ�0B4 ��¾.���Z4��G?ҖtC����׆��D���i�Y�e�6�/������ð�1T������#G�G�0�Hנ�# ӔԮo�oG��7a�{:�T:�����9��$��M���^�m
{�~���b@�����<0�'�r	������n,�����7�;�ݍ?��"��9:X�R1� Me�.�,�R ����!}!*��^W5zB^�RB`�r���\NQr���&�6��/�'�}�u5\�c^D�t7#��P`zˡ�%4����p̣�'�2t���N���f#2qR_'�ƛol�S�«����;L�䍚(�h��O�1u�T�r��x n�2bK����n2NO�)��2��]']��+���Ε�R��۴2Ϳ-�L����g�h�#�L3n/GU��x[����oa�2|�[����ϛ�ġ�.�G����f�nX<f��,�_�W�=�[����:
�c%��H�e���U��TE�X�p�6���J��*mD�~V�\2is�9���ϨQN�{��YΥ*r~����Y�Te��(����/�C^	��*���+�cPw�SY��/އ�Ʒs|��b/\��1��7��i/������s蚂�ZD}MttP�[p�#>��b�1n��iS��Q":gN1����l<FLT�j(*�ʃ����6d�����R9��I�zq�m5x�߇�5�`(+	H���?h���܃=WH�SR"K�wei@2{ Ew��������4��� �z�r��X�\�7��P��0�yI��O��`��q�K�k��5�m�q�kv�<��y~7ml���-m�#��,�p�����C���Ç"q,_R���81��儬��]W"5�rv�$�Զ��#R�>w.�)Ǳd���@`���y�ĸw6Ǒ�N���;�"�i�j�a��*�plk��{Z�|N9VR���M��ה��d!���i�o�l[�5�#w��3q��P|��S|���j��q=fNϧy�q�
+V�����w�p6%�:3:
�*��2�\:0x���{��T���b|��7no��7J��(�ó�j%�_x}���������5���kh����^��Ϟ�%�K0��.�b෯���kPR��/_�T2��u˨P5ݏ��y���_?s�y'��:�޿ �y�Uy�,<��:y�x\H�[{���B<z�<� �Z���5���)~<r�\<��6EmA�uI�V����?}�F���;N�3o���kN�@[� ��L���������@�l��%�Ȕ 
)��gL��<�����:p5������+���#g���)m]�CXD>b��)���b�Ԧ�E`������jƬ��6�؟���PT�o!�h�$3�v_ɇ�uؤ����y�/ _9%@��'�g�`�_`�+��m�m�h~c�4n	ǂ+�IA	�f��ɹ�'������4�l	&#>Ի,��;�U��`�������#+�N�aӮ��bS�rY1�;?o��p������X�7F ��i���s��;�Y�!��,�a�t�!�6v�d�?^{����v�[ 	��m�l%�G����	��\+��mn�>�l��a�	t������X�t���Zۃ��Y+%%8,�z����K����&d2��I��dY�Q�r��#ܾ����M�>d0��Zq����F�������
�USf��PU^ �v��Vɤۮ��~�$�@>0;K6Q'[���T��+����hEiQ@FzX�I�(��Qo���7�������E�����?Տy�S0��X����
S$���F�?�&�d������X!�VO`��FuyiR�<#�)���C~� ��}���c2 P/�	e{���[���H��B;oH���Jں�d4�S�H<ž#�h8�Ѓ��ݲ�c��e�鑼C��l������Q�x������Kec+�h�R6�9�&�Y��퐟9l1�O�qlj>�3����#s�>�&�ە�#J�f��&{�j�;�5������;�G6�{��zEu�T�����L�'2ַöQ�Re~b�T�R�i�pD�v��4�2�0e>!%M�y��X��8�?��LeI���
�/�F���1�t���s��˴} }J�*ι8*��T�g�?(:_�8 9����2� ��D�r���I�(V����
{6�ux�8�3d�o�y��1�e
ѴH?�w�CKd�|-�Ɣ>�Χ���G�J��s9�\���q�1u��2�Zv�g�I7SL�2N�<�};�b??��g�9�d<I�'O�����sL|>�_P��0ׅ�)M���=# %hZ��6�3���/�D$����SNӻ����my�4b�]tůfN��o&���P�%�����i�g����х���-MF@"�H�E�M��K~�7m{�@�Ӟ���|��CCCC���ԷN������P��U����N�1��I�E����n�1��þ��<&^#她Q@(11]~�-}�w�HA����^T�R�0�%E�4Û���3�C��k�����dc�]5��FKsy�/���ϓ��V`��� qß���`nN����?�%!/��W���DZ�d<���>*%p��'Z,�C��=&�]!�qw���P.���<A#��w�G=Jr��F}��o��xBؙ����1/:8s���:Ge�԰(T�gpyЊD�� j�?�Q	�E�	�[=�|1�*w$*�a�r���q�V*�PY29i|D�.1��烰�y�������r��e��"�f0��bv���KAK����r��``Y    IEND�B`�PK   {c�X�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   �m\X��>}��  .�  /   images/8ddf307d-15d9-469f-99e7-c830f4f75d99.png��W����P("MJ�zA�4K�/ ��AJTZ��*`T@��.�I�MD���v������ι���?0�1�H�Zs������RWG����Q��S��� �r��0��=G`}5ePI/�
��(���7��p�<�
|�Q����J�X^W�2`v�una�R 	q;���Cb�_mcs_�#�XDz��̡����JFI�{��6��LtN�O|�oz�\��xec\�۾��_V������~��ϗ�/�0S*`=8��?$��b��H�9Þ]{A���R�����i����Q(�{����i7��}�9J��.��7�<�����N8��?FQ��z�Nb |S�?���� <�?�@��� ���;lW���'�ׯ@'�SB��g�(�����G�fz ����^�t��c=*!��(�xa��?F������A��ZЌ��y�0�VƳ��Ê�XH���y�F{^5��B���t\9�?��]��8m0��m�sU4�y���׽F���B�����1S^:o�:Ӏf5=��V����h�@�>j��L�D�lQ��K��F���Û�_������8��d:��UG܊��z�?�ۍ��J�|��T8ʮv|\8l��tRѻy�9�%�&ߪ�q���쫛�9���k0H��R��E���"�PG�W�dt����	��Ovi|7;<Yv �Rr�)G���HB����V=�tlRw��'���j���wc�xh	��QR&+��I�W��9J��C�'�.M�
I5Y��Q�s+o�D[D�"5y��.����y�����{�<<5Y�ƭu�WD#�x=�N^Z��{vR��dܢ����%k����3�后����=��ګ��L)K����{��q�Z7�D(�#��P��
h�X='�,"�8�={=p	�=ł1-�t��1Ũr@�a���"ZL-1�����'+��On�YH�Bsl�d����t�6'ܔ�nC;D�M_��j����ՂVd�R�3��9����J�a��X����_[eɰ�/J5�����0�6�V��Le2�,w�
�W�������%f�<���t���ԏ?\�V�ԸE+�B�K�39�����ɓs>���!d�>~DE*���P����Y�.?�6�X99��}��O\塽lF��������5�u�Y�p��*R��QiE��i9V���]Pk6���ጎLj�荍����7N��b́b�=Y)�I����]
?���D��0�k*b�����n��f�|#�j�ӷ����4�"����&w't/�ZL:V�'}2���	���2J��5߻Br�qz�?/�<�	B��X]c��Ȭ� f��������ϴ>��>���W�γ���̟��
m�ϐ'%'�_����ܢ��Ҋ��lj��_���
�+��	nWw9������'k����u_�s��u�S��0�ޚܐ`�ecC/�2e�/��1�`A��9D�'.xt-h|�mٛ���*��]��D�)p¨��o�z���|��H��0�b�!:�٪�=��`� gt�"%%���-t�����=a�сi�;&�Hj�~�)j�A��r�+���
1E�i��>
��{�I�v �J-���ѴN��0)w�c MJ�3GBHde�׫�'jY�>�>j��9(r@]5�A�+�ܹd7�wo��K\���n�R��Y��׉Ӓm����Xz�����+����No��i��-�ʸg�pn��39�G�vNb9�3����%鹆]����5_��zz��_"�|�n���5���Ժ(�Y�&#��N�`AL?��	��̞'f�a�����!����5����:q����A����y�]&���g>)Q^#�ev
���4Yy�a_q\bg����}�p���֊�)*o^IV�D���mȉ���}�.`B�A�N��s��dd�`�h��eiG��a��a�1?����ފO��V����k���nq	ݶ���M���-�{�?��������;��[�Yad/�h zC�P��m��.伻t��ʟ��J�����?�NZ\�`F�<.&Ls��el��w��fT�mP�Ϟ>3:V�����F�DYM/;���+�6c^�(Di���{�
��k4]�(��]�K%#fb�R}����E�K�k�i%ߪ@T^Ŭx���mԃ�x
����^��$�]��7�G�G���h���Ha�ٕ8}�&����v����2X�-��W����� )0�nB��p����"1E|KB�$�Y@쮩3Cx�$��s���h3=���=N��cl�ף��0�@4�m-W "ܗnaVv���&-d�5��<��Ä����
m~����vŃ����>�>�-~���$��vСt
�wC�T�����J-��p�ɸ<�Ʊ�	���u���s
{�b�}���?>�e���Hl`���Ւ�b\�_�*o�XK�@�8f�G#>A
�/�
fO���[�I����dI�+�GF��e���O~*����bT�?oV�/L?��w.�B?��3����n�7�]�	� U�w���κ�p�L�^1_��LŶ�j`h	LA�Sa����r�*��*3~N��rQ���w��\���=# 4���(�P3iQ��k"��t�G:DL]Ie��F�S���,Ϯ��D��/�3�[��J��6�oRғb��#��*�?=�r�����3��y*��z�ҧ�/����d�sXq�d�vy�y�j̶�Į��qXm�r�����[��I XD	c;w�����Sl��#�s��~|$�����'�֯he&�'*��7�<�:x_��ʭ�f��P-����9i�y�}�w��^�U�_��FHno����.Q}���i��t8Ќ�5��B3/��_\�Ҝ�!-rvs;�f��U����ֳ�����,!Pz���R�ɷ��ӹ�Yﶾ�T��2Ի�ۡ}v<�E�d�m�S��x�Z3ÑΒ�ӬI�@Z���1na�LpZq����_X\�W
$�u�B*����!���������#:���a������sN�j;�6	��@�D�0�,%t���_,(�|�UV���*�`c�-���{Z��k!Q���_��A��p@���G2X�)�ՁQaf�=I��ԫ�qT��,4�X��x���/QcqFvz�/Ց���*&7u�J�F����S�����C�V+�w�2��~�����fΟ~��K}��	�8AC�ݸ��}�ԍ�a�[X)J���J�	]�K�\���_�?aX�߹>��qMHtÌ��[�12��	���Es���@$&�S�%��M a
Q�îo5(A������5��?<�I�K��@�<^����Xφ97����WxJ�Is.߾���B��R�[:��&m�=�/��{1C�eoQ�ޓ���x1̊{�]����2x��Y9X?����TE�'cy/Jn�6K,�T_,^t�=ɷs�[{��F�KШLy��{?ȵE[�d>h��舡��N1ej�����X������m����L��L�FP]�Nɩ#��9#�W�ڿ��1��%5���x�[�I����_��jl� fזħ@�[���\�l����>�z٪!���Y'
2�2�����O����up��K������]
���2ͷ�c d����֖n[�]��C9;%�ߋ����O��bǮ�m.z��::�*�3p�ܤP��ϖ>U$�����?��c+���1�5���|����4���T����sx�;X�a�2����m��)谺VTW�Jz_���f����&[�KHE���T��;f��Rse�aE�2ݜ���B1À`�b;@� @S��Pr7{�~xL����_C6q�acǯ.�ĥǈ�ό�P�|+�D�x{#��&(�~���{cB{8��s���B�$�1t��R�mΓ:5(��z��˥����/e���RģV8���e[���|L(8"t�����U��)�,�8ݶ��ۍ��%T��_��z8�	�a�Y|�q.R*��t>ޯz[�'�!�%�������\���}��?��5�]PD�xҺk&)�-��7��R�^������~��$�G�.�0���g��4��R@��[^@�o���v�E����������6j��5����NW�do���N5%�<��JR/��Kk�ؽ3d�;XzT���J�
�~#b�=��HxV	/���i�m��)p{K�
#�N�ǥbn��L�����w0X��s��#���M��G�����h��#�M�o����*D+�R�>CŰM�'���|���>N�4Y��y�a(��/���۾&�MR�C��[ɫջ�?��Z �E:Qb������Gjڹ	'���k���!k�}ٲL~���pXr?�l\x��z�Y>�ܱ+�z�
/r�D>O/�ѧ�ge�\������76ޅ�B55rߐF���d�j�p5D5�D\�|��B���s��4L��T�z_t�g}xM�P�~��K����� 4�W�z��7Ma���d�k5����(-��� �ο8�X#Ďx�|m8&w���dȹ�#g�V���6��~]��xTw�C|�]Go7ojW���5��Շ[=���
�I��j��b^1��˥)v�a���{��>xe}�ל|]e#6�	)��b�{-\��{i��0�"�g�t��8�O�X�l�d��ޝ��YҴ���kIJ��Í���]D�c���Pnx�0n��w��9�|~�%�+���K��>)	OW�zS`�.*x!�;�T�t��A�4�bK�$R3)�kx��ߚf$ػ�L�P�2[(K��J��5+��$a����m=���=t�8�z�5��x���#���f}�b��H{t��%tm���kB��qS���}���Nݲ�s�XҾ�3�-	�PO԰��>{X��P��;��tr+n��EG�O{niВ��@�{6bsd����%}lmtR��K�FR�M�c�����D�{'��n46�;�(�Dl���mE�!R@<�;�����L�H�oT�&$�u[���bf������!������"��j�5=xU�E���9����gf�d���waK�^7�v��l/����Ǖh:�h���"ƶ�r�"6z����I`R �?�}AS�Eb�+��δ��a����A�+o#R9A��GԲɂ�d��s��Ի���>3��-�Wi���Ա
m��ݖ	�I}<"y����߹��k4��e䖵�}�+��cR��2A34H�H9u� �����4Z���Cb�3:�������)��篾�Tc�7�D��A���sqd8�@�����85^'�wl��|;����*
`��B:�h�u��k��^G�J�|Z�j��Z4�)3��+UWoH׏����№(��äݧ�
��!�QCP������o�9R����w�JWW�L�R�����Ċ8."�NK�K� �¥���N0w���� Ts��8�><T��Du��p٭���m��8{�I�Wd�/_���ِ��k}]�Y���|���s�����S��8�^(f��R�?Ft�����ړ��z��f��PVk��a_���}0����������e5�&� �q88�b��ڤv���I�md��&��H�[���3��/���P�}�L��D�.�y�SI��;H�Ay��Y��*��L���g��^ǭI��oݔ�_��mqB�*�K/rїϞ�R:F��7ż`�Q�W�#�t�%�q*��xI���m7�q-�w�Qr����V�{����bo��']�d/F\���syn�B(6���JQ�/k�Ӷ �r�dF��a�;�`k�t"���y��hD������2�� �����l6� )�VbdB�RP�./�u��«�oV%�T��55�k�F���^}2O�}��V�o�[O� 2C�����"�<,1R%�����>ju�tyh���Y��nw�֘KfP������.��6㇆�Hm���_Z?�i��5J��A�`&�pr�.i� ��)
�~f����P��v	]�gJp����G��'ι�A��k�����"2.G<�D�ob�*�7h�g�"K��f&��r����ۦ�M�.��Ó�����[}kp�+A�2%1g�9|�X���r�e��H��AG|ԩd08 O�i����}:���!���'�����cr�j�������KV�O�6>-W�wn�\�>Wc��h>�
�r�z�) n��4�m���^+��Q��OE���([c�T
�;�[��X
'=_	AH\dF���#�L�(M9�%��t�5��ʍG��f���~�G�,���b��~�y\����-W�����pf�����|s����bp�:���o��u�+��Ii���қ�Z�"/|?
%/�����R`,�>��2�.c0��jĘ���Fj�ώ'�-���O��y2M�o���	r����9%�?�QfEJ�1�NU3_���8��X�Ђ�8���o$�%0��S�3����Z��v9����d�����+H��2���
S ��9�8E����G�ݭnk��ψ/l�c��,�7��"'��oe�J��d��2�~��Ű��;�A�]�:^���@L;�S��%�;���p+;ӏ���P�*�L!�A9̥I���hU�T��S�3B~���s��d���F%7X`���=��q�}R��4��Q����*&%�Ȁg�t2eT��M�≾&���*dJy�L����T<�ur��qb�o:�7�-}2���O��Vz~,ZMÿ<Uaԑ���%J5����*�$��E�ꍇ2��D�L�4��j�S��&8v9�8�R!UN����+�ʫy/�d�ߎ�5�bd.�m~�e���=�la�h�i�FU���A������JJW�w�KG�~��O'WnT'x��'�&""vl8̿W��:�v�x����P"�9�c2����B�$B��>�qwV��k���鍺��W��>����ɗ���(��h즮H�b�?�^H;�{̢v���t��Pc'M��&��GV?H['�~�J�X�9�f��H@D�(ڳ���_�'�9uJS�J��d��xcA%��(YP���6]?<bQ&��o�5<�.(�^7��w�����Z9�t�Q2-�Q�ac�|-<�o9"n/������L����^ڑ[���O�����o.�Z�C���F@�2��1�hV?�����*�?�@H�%�싞 ������q0R�;xz� �|�ۏ�G�*_kpz=����އ]�� v��b�"|ˀ���f��6)�p�9$��g-+�>�~��Lbƃ�IX;�:i�����/r��̼�1���߽��"�_�=1mZ������T��,֢�ȗl�B�5(Dc��L:r��jln�>��O�i�4Ji�J�W/ �{s�����9}��"�R�����^�LG�4A,����ҥ�0{�����Ȥ;,QC�����Kj����6s'j��j��.�qH��
=���Rz�X^򕫞�t��-�ρ�}�Ӧ|�Y%h��y��y�LV�rB�q�n/%^}�Pp��ܦ�߆�M#"���;bXeuq�'H��3���a~�0�2=�Bn�m
�EvQ	��>��Iu?~��Pҿ��S$o�П��O��1|�W��%!}w�ǿu�Q�7�۹4gLջ��]M�#<�%�W:�
eI�~���=�{�?N��1�l�:a��h���)����.n�-f�T��-��,;���8�Q�
j �Kiz۾�i8!�3�/��T)�����$�UU	4A]&�Ls�i� ��\���\b�e�*�K`4�:��c�����}EP���ǳ��-�:���������o����Z�R罖+	��/�n�ܽ�D�:~.���'��V�G�/�s�d�7�il/�=&���(�S�n���}\��h�g�����b���`^�i���t� ��2u313��P�t�\��E�f6�hIB���sC	��/y���O����3Z�l�ʉ�����Gjg���h�\͸�L���a�����}y���|\�KQ��	�����K�&�^�vO^:1��ELXn|�FAF�2+w;*pR�?<�V�����!��s����j�I8�2
o�i�֒���r+7h����FF/+{:�#��N�̓�7^ȊS��J���m�6�% T2��]�1+�I I�*L�	QH!%%�}��nQ��
�������/x�wV�9���i�|�(�*���I-�>廝�8����%g�cA̩�����
�y��(
��P &�����Ƶ�>�D��YS��;#�,I)��s�{qS8��P9Lqi��Ue%y��)Q;��68s��"�Ŝ�U���$��!���r�;�ԛ�o9�ǁ�p2U3���!ۈ?��ۋ;��ݺRr���50�eN,���o��ܡ�¢�6���A������(���,a*`������Ʀ?k���x��u�)�ZSr2����y�����7�b�d��}E�JӃ�AB�Ҳ̗��h��� ��'��1���F�|?�֐=�Y"H��ۈ �@L���0�Q��cQ*u�0��A��l	�O%'�n�1�1K��/C) �
�ȱ�����i�^FX�KtO�@���E�X��D
��e�&H �'Ե���7˚{�hpŶ��)c�<VP�Cr-�>b��Q��F1g��?�kek+�"+6�@�~|�˷]�ܿH�[�y�^�Yj7첾d��QJ*>��,��k=]%�N�
���+������P���yK��jQAA�m�FA*`[���|�x���j�lέ��v�T$*A�J�B��o�����vK��ӧB������E';�>H�.O��q T�i�T���?D%�[)���]�./걇'�� Lc_!�W��E
s��Y-�DuG@�';�8�c`qb�:X�/�����̒|%�'�/��0JJҚŷO�o�޲S���pi&-��O�������(h܅���ޅU^�����mh���Q���+�,n�q>9�KF�)��<>�,e`��a��OQi�}C4�	%�y|�`�%@���
���<���V�4�,����</ā�ԯ�=��N��j��{��͆!_w�F���@)��'7�/ב�Ar�q'�B�\�̲�yu+��+�`S��NJ��_x�����(�����l��9W}M��%O�`_����Z�׎��m�x `ݵR�Kߧp��ɢ�<2q<��Nl�o�~ӸE/.�[�ҍ;�[<�e�9�m����F�8"�EQ�R�%MV��e�$���)Hrٝ��[�hf��,c�7z����,��U2W�q2�i�����-4�v�G.���pZ��P_r?���?�Vs����m������}=��i�� )�~IF$��=?H\�h���0���C���
N0q��K�6n�7�G�g�e���fr�&���F<��3��f�ؘ=2zy����Q4�),�%W�SVo�n�����K����k�^x<��ߏ$�أ�_���(���??e�����
���פ�j�R�-�Y,��[�Ck%#�to����[�-�VB���W
;+�v#M�?|�շ��-)���L*�%'�@,�ΰ�n{�ڢ�cV�{�⫉Oψ�7�S3Au���sC���lzb��Df{ǉ$"{*@�,�?���UL�>��=�,�)A����B�}��Phwl��"��VK�
Q$�P�Vtp)CT�B�Р��Mks�{�9��:H4n��>I�������*�̢��6*��#�/�(�3=Z�d��3f�~�.[t{L�Ȏ^�j?�ƥ�Ų���N��c�J�Q���4%�neȳb
�M��$�ώF����.Ց�ڠ��чR��Rs��l  1#�H�ֈ̰�?i����A�׵i������"d�Y �NѮa�Z�-��q�������%�u�� �
"��-t�>���`�g6�8�6�Xu���r�a����F�_&x����l�(�`��ђ(1�h�f�ba5S�1�=+����r	�AC�e�>�>��9�$(K����П�W�l0��Ax��=W�Aͤ��o�,�/��eG�:���U��%�d<�c�tu�qUy�|߃0���a:<���ho�~��'-�l��$��V���Xe��i5�1R!�u���>wT�L/���K���������'�-��,�=�:[�UEh赈S)/������v?$�V�.�}Y�|�v���3hB�ݐ��r_�ο�����gM�%-'+s}������%������N� ���<�N�<~l��C����������dt����|B$���RK^Ϭ�#P*�D������ ���.��7 �#9R�A d��4)�s�t�(��T���T�uw���!�g��c�^srb���o,c����2�3���Z%֋y@f��J_�P�`Y7���jd,:����sx�m6ĥ9u?IpCe!�4��ha1)�Qp�wl\��w�x�Sh71F0zX� C*]\�g�ؓU2?�!��+/���7�������#۟���/{_�4�"����V�Ć%�xx{�[�v����f��aM���L��'��;��"���s��p#�}v�҉�y�2t���b�N�c����8����ԟ��'� \Q���ׅ<��̎��"�AO!	(BD��)�6��@�f�>B�!�$)o[��+��s�]w��D:{��l�f�"��Zc�����8@͔!un�l�&#����R=���aL�	&�l���������>�K)L�p����\|��#��J�ݭD��4l���`/#�h�i��A�t0Ec�Ē��$\��m���A��5dcG���ߢ��i��|B�޹���)����2���|�����$��m�<�lɞ��ؠ�br���~F1�p�Y�����3��		ckC�n &�)ߤ��� �@D��� |P�!�������1��sy���p�S�T���N�Pн�i��q�{���	Y���D(m��e�1��y �hͰ���о���iG�j�8y|���[�8�J�:"�Gؾ��!qK~�E6�Q;[h��Mn����%H��KĖ���LV��L�s�;��w�� OW;�e�
�0D����gr�I�	�^6&7�1(h��(1l+�q���.�(�*�Hq�p)|�^Ds��O��%gj�R�j/\jL�W����|�'����ήU:�l��}O�	*�U�N#{�����F$u�قuӊ��M���_�O0f}'<�b��T ac��&8�>U���^<�X���ԗ�G���6@Gf� (���N��Ƌ�=�>YYN�)2�k�LO�2����爤n��cALjD�R�4@�)\�5yF,2rj�3���^��vy���\!l3:�P�w���CyXvs�i�+!��i�~��7Tq(�,�����/���Ċ�m��@���=���hךgG�`Ǹ�Y�==N+]��K�!v�lh���F��;����O������c��z��u����#�'IK�rbC�߰�����Ǽt;	=5$�O%��.ߕ���㍧�rpv��)��g�,�O;t����<n�m�.6�tv��6�o<����✈�~����Ǎ��e���{/m4m���cN��d�A���Ȇ��i��}�J[�<�H�j�Q�D��^NA�u�F j�%)�_�p�����+xU��^�V�ͯj(�UPM���
�[bj&��A}�v�ݕ�7�Iܭ{xq�G%܆��)�>��F�C�A��7ֲ.��`�N[�����+�V��c���Anp�WtQ��0vh�NJ/G�nx�Vpu���&<j}&k���2����~s�0-��|�F�����AX���td6)fɽ���"�"�?O,¤o�m�@h�R:/�[�|�0`�F;��b(Kb���(�6xgV����Qil�bHܗ]��F���.�PI!�M9��¨�,��),$�X�����a��t�D�xNVu�|-D������!Ww��&}L �<�b��$0g�����Bd���6Q�\ZTv�*>�Ȥ���J�ޕBC�jѐ�)R�^�� 3~ك��ڂ�hO����h����T�V���6�c:�^�h4�U�s~�-�	���sh��u�E�hH��B��p��n��Xa�H���ι�_�n�<cQ��I��RDC�*S��^�Wi9),�t��b����R"��.}xa�'��|�FP�,���?~���3�<]�~R�N��"j����0�#d����~�|k9�q=������u���9�C��>v�h�������7���ߢ�
Q'U8hG�& ��%o"�B���B��k��W����^�~у�
�b�#a�/�KYa,�:���Ґ����&�$-�*�=����̶Ƹ\E>�~4�ǭ"�$�>�Ge��e"��h��LU���IԸ�I�Yax�~���aL��%��R�񅅅�i-�g(0+5�a�8G�=%d���.N% �9���������>Q~��,���x� �W ����6'��ym�Ĺ�ȼ���FZ��j:K���h]��ޞ��o���63�۩��4����#��K~�HEo<w��Srlx���e��$p�2�3�t�mC�mc[bTlV�Q�,ibw����|A5P� ����l�ٶ��]Ȃ�`�Ykaa�}�.�7m�����C(c��J�y(y���A��9*�v<������{cayA^�Q�-9��#ד�A �JԘM��)��!�Uu�-�fNz��v)��]�+lo��@_����;k\>��.F��r��|t9Lά�<#K��#ǃ�b�g@xCEocn�HS2EK��}r��r�����,�Hɤ��:�L�m�S�7�� O��4�C��_>y�60$���y�/�V�D���s�#�m�<j�����yJs����`�E֣�	xe\&�{wIq�a�6j�"_�˝q�����=8��cP��?��$t1�m�_�R�ALR�GG�u�k����Ͳg-�~��u �k���e�$�=\8���ȩY�̡���q$�Xc����.��o��|��oUE���\�J�B>X������H�g��:�(�Gi���}��.~�d���Q<�v	�ZR�_6��CB.�<�b�d.����<fnR�a�:Y���k��c�Ln��@ӿr�"��������~��k�҄|��8Z�YD�Lh�]���� y�W�}��~Y>���:D�1�gFID�)��)O�C-�n�ͻ�}���A��A0��N���L ��.6���K���ke�E�z7ZOtL�S�����֯3$�IA�=�މ&�R�A�|��Q���m�i��i�@��w����G�jY���Z���$� E1�Zl�h��._Ω��q��q���Pݷ0`fU��k�2P�������\,,����F�ZuN�@����GZ��Z�L&�A�l��f��1�v3�G�QD.�%��A��I�Ă��2:X����B�%�߈eK�ߘ�Ԝ����7�%kyh-�]�k�O�]�����ױZ�U4���ˁ\� ��>-��6��E��[��N"B穒�{7=.~�'���˝����P��a��>���M\6����ۯ����MB �sS�6؝\'f[SI?�����%<m��7ޓf�^��`�~���Q��U�?�1�$�Ǧ?��Z�K�U|N$����Od7�L��;:��#�6x��ֿ��6�H��N<�q��{�c�jG�w_��?-fP��b����2���܉.��bS{�x���l�ɷg��$�u��¿D7��D�����n���:M&���2E�̞����Dy^����h0����:mp5���9�|�k��\��������KQ"�F�����_X���|��7�C��dU;d,�i|��
��\�/+�'j,�I����� '�,s=� B�v��/�3k߂���0�c��X�Fe�1�#�N���s�(-�J���U�p���V��l�v6���*R�N�Y��~���˕��"~�R������H���q9�f�`'/�V���l�������E�G�d/I����ᇞ���p������#^��DR$P!�]3��Y����k�y[�RFX�.
D��cZ8�n���Ƚ�)����'PW#�e
�F;GH�/f|N�wgMyb&���*�Gp�}>����2BH	Kh���s����Ў�%M.
ț���N[�/Z��͏��X��/�����T�nZ1��_E�����2��q07���V�����˪���VL�7'I?I֦|��G1���k���uk$�,�WT|��#f�D��Ԓ��cN��ڳ��Ye)2��_���k�%�5�n��2��*L�:*������v��3ҎokJ�:�	2(��ʷ�D=�xt��Y��I��8"gX����&�f
��T͊��$[ƚ��>M�bB�0g���7)*Z�\ʍۡ�2�9탲��l���y�����j���|�k�z����;���Q��������ȿ�*]c���}��:sqK�o�)h�]��8�,5pE�츏��˅�C~󆍀��s��M+u�{�4��7�~���
��m1܈�ԜI�>���_�P7X{7�~f�L5��q�|u蠫[�uvY�E&�M�wl��;������Շ ��ɰkܳ��w�b�S�(y{����6����!����'k�Ġ�D�6)��x�����*����,!F6�AE-���+�:.��'��2��)2�1�ӿ����X��)v�8IQ�uU�}]���ov{&p��4���o;kk������)9p� �����XkV٧��������cAGet�F|����y?�#�����~��-㦢9�vg*R�Ϲ�~�pM�zA�7x���ȫ�Y��w%9�����a�����&8����$h�ѝ#oaă ��,�L#`��Pb�7q���v���e���G_�����k�z���$*�+ac�M?�	ђ @�s��&Ǡ���ۘ,]j$K����ȥrw<�d�C�>j����^B�r���SX�WS�����g�^ۧꝩ�B�#��V͟�o<�viX.�;���>�� Za=�����bS��e����X�g��.�;��?��?��3��Pq~���l"�<��iBD�c��C�������Y4^�o7p-<n��@/š��Fͷ�2/�=;i��L�oϩ"*T#Ya &b�u��e"W�����X��A�Ǽ��4G�FҚ��dȥyq\G��ʲ�ԃ�E�&�`&���I��Qe�cY t�iiA��U�����s.KG"=�3W�
4}������B�MBx_M��L�>/�q=sP����
��F~P��Wl�N{��k�֔��]��,bAk��M>��M��[k��ח���O_���M<��K�Ɉ�����X�o<s�KH_�ç�R��z�����^���w=��r�t������` Z5Ԕ�
8�]+�����:p	r�j$�S�
!��ܑSRj��� ����JuK����a��cb�T���}��?�,��x~�]X�)@F �����&6k�;�?��ޚ �Z7vj&o��"bS�%��;�I�gdq�rx2H�"��h��}zٹz�X-S��y�Ӥj�F������l�aӫi��J��P9-�]r����t�w��N�ϋ��j�4��^K�����'.i(�f�,��L�Z�@q���o��뤲��y��mɠI<&C�x_B�.d>[�\�ar?� G�ڜ�f�-yaR�{�`��ܐx�UG��OΓ�Z�GMC�C�s��x�[ܷ�7���bޮ ����:xJD���ϱ�,�v��\@�ӨW�ID��B���)ݡ�8����Ã��#�٣��R�Jb�<�}noL9U�.��>��y�}c8�M������nZ	�7l�\,<kߪ���o��6ʊ}�0�aCt��X�!�Ek�=0�9�M2���;���|�u��,žjܪ,|h�=�)5I�����?�Bفr�;�b��a��!^�I�I���L$�?d�ؖ����G��X�K��u|�c ����'��!��J�.�AFl_��y����&>[�L�br��j��d�@��5'���A�m'd�ݣ>5H��L=�(�;��=۶<��k�̌����Q�&�ݕ�êM��;`�ah��;.���ˋ���?׏�b�\$�8�ʊɍ,�q���%�oP�A���d#��wk�$���������,�]��i?�d��>�_���o"PUu��U�>|���Vs�K�a��%[�Q9t]���D�ʏ{u`�uE��(��Ld�>��A��GSeJ���z�)<1T�$��y���~����%��e�$N���z��!Q���L(�%�2��/��6�L:��ٜU�4�`{y����z�o��f_��r�PƩ�������p��5bE�6z�_����&,����Q�v2��qɜ;y������O�\ �e��n�w�67>����ȵ���L�e�%LD��?rÿV\���v�.�j�#*�4��} �����ۛj$V��d>YjiI��7�sF�)C��@�xuE�����c\�k岙��WH�o�(�UIɃl�t�x.���*0ټ�α����h�����|Y�C.bi�]\�� �y����i��C~#�A,0��*����)S�	Ќ{ݷ̞ս�++�6q��+c�D<��~3���\$��l<j�m)���g�Y^���0�y ��^�y���ёM���_��OZ$�fx�nI�?Q[juF=T:]��ĩ��7H#H� 
�\ZþԶ�I9W�mP�K��Ё�O�?�G���Cv�4�mAM*@��E�u�⟋
)5P���7A &��C�[�Eս���H7�R8t�tKw���]C
H� -%50�H�t�H�;��?��2�c��u_���v�A~;w&\�%mHQ�}풣���}&��g���S"A�P�����:$���u98/5<a�4�Р�/��`�H;���0 X��x&���:E0`�-�a��v\yh�K�����7;�v����7"���Kd����|8]�ē��O�'�7ʴ%j�ꪧ�o6��ie�b�x��	4ks��d�Z�����!����Q�_&��*��$�9�`~��j��¼����Z�
]�P���[غ1�_D��&����@6��&w�B ��ΰ:�a%֋h�W,͉
�x��vp��> ��S��d����5���x,���l�ֲ�EG_ȼ�A�Ǟ����,����2� ɚ��e���3Ĩ�n6���z
�ښC�,[Ę�&�?%���Ц쮰�N*��i����G����J��?��E[�]7�$'�7][F-D����S�.V��������V����p��C�]9-av� Q�U�n��_�|<Cl8a;�iϔ&8�8�r%	0��&�_*�lP�}Jbz��O9Ԋ\©+�J&_���y0�B�]�*[��cQ�8t
*���� �s�v~'Ӷ��w��P x�L��L[�b<	��z
Nr3��1^�b��B;��R}s��F���u-%�M��)<��?��Hg�>��H�N���ZTx�W�a��~�P(s�1� �R���*#�e���~$����G���fh1GOn��&�7�um��2�vA���,���ϛhG�r�ؚO=�a�k�L��y�����)$'GP�y+H4�-��Lڠ�LE2��6wN�~��UTvTt�}���dX�ʒg^��������uk���?��f�^�ی�&�;0�YC�?��f>���5!���sω4��6  ��܄V�����>`�Su�*�w�R�䳲 ���O�fzhO(�_�O�!�ceR��u>���.Ngp�hb����1���w�OB�ۊd�����G��4��ߊӞ<nl��m��9�Q>1H�֥��,�Wn�O��r��Z��2�rC��;�ǣ�����kw��ٶ4��8`��XjfHJ*��&3��Z���໡b�Hn��Œna�fq��4�n�[]�d^�ӣx%�A�8m�09i�����/��8�9��S"5-f�b�N�VE�{WT��)*K�sH�gO
�p������� m��^!(���O�BMU���+=�ʃ�����y+��JFw��^�)TnO�T��l3{�[z��H)�6a���j��$Dт�p���Nv��@�d��`"3�e�B�<Co�����fJO�E����\{ؐ�
a����G�tk��G-p�ۧ������e�@r�����ޟ������0����]_lD�~�ih�R�3��D��t��!�eP��k��+ퟱ�����ul�/@�P������������5Zx�z
�oSH���J:~��~uT�*���w�:������QW��� ��ӌI��ɦ��wPI���3g��� ��Ѥ'sm��w5�(�Ko�|�e���1.�k0�d�[3;o�����ъp6�yd 1�V�tV,�
��܌�A$7_J08�͝�����w�M����1I��n�5����Oȵ�d��+_�q���l<H}U��]M����MN��A�vݯ#M���r��z6����]�!��mB̈��}�ߗqڏo�^i�GKf+���5�W���vܒ�H-*9��A�L�X�����t'�w�3�S�%���J���C�4 ���WOP�X�Sa95M�,�sp��R��"iy^(K [��=��V�J��A��L8f�3����K����ݤ�A�q�����k��sЊÔcM�9a��|WΨj�F��M��������1U���L�j�&��A��'}Os��d/@�\S{3��pW��B2���.f��~$k�^�����{̏�&ĔV:F0mX��/���k������z�瑾�/�${���S@�����7�6��X�Qŝ|;���P�d�-J[��!w~�<3Sv�Q�˥� hg-�:������7�'�f�!��\���p�ĜB���9=f�7��D��%��{����#/�|;�.O�8A��~}���Q�P�d�%'0�j3�ɗ�qR�L$Ϡ������y|J.<H��ܰ��Ӟ�շ���=}a�g����amy����Ԫ,i%y�^�,y����uOr)�z~u6��o��4��x�R?`yv���9���.��x��*��(��` �iV�RV=>��Zd����f0E��*c��o����D���G�
!���<�A��U������%Ŏ���+�W�(�[O���~�\�|[��L���=ƌ=u9�eA��v�<N�o����	e_	wI��P~�9*��C���oͷ�b�࿃�8d:��)�h���L��	��w?^�!醞v+?�}��Ab|�H�1��%ǔz=����_>@���`D/�}t�G!��	��y������TÄ�S�f�� e��k�_��߾;�@�aJm��s������vS#V6��l��V����D�`��%�� M�>v�=
���Hb���ӹ��y�'?�4)����7�eD
�<���t������0ǂdp�w��~�fJ�87,E��xr:vƙ�Co��.<XY�$O��4X:Xs,hr�/;݄E}n����]�R�G.��먌`g�>`��sB��^�*���/��͎�Q�W9puCh�F������' "�X�!�p��<�z��79�0dP�D�]p=X3�w�)���9)�n�d�Va?|+U+w�b�~��DI￲2����dԬ�V7�=�7�:߬��C����|'~g*{�� �ߒ����͓�#�J8QK�ă`�g�Ďo��b����O���a���.}z;��(��a���xy1kA�{��3�~_jA���xE��L���ї28�]�/��QF
�^Q�6�Xxf2��ɪx���F��4�̄�%j�K�k;8�%j-N��nr�ҽDv� IU�*�y�D��o�Õ 
J��Qz��hH�o�\�^�N�]��U2���F3��ؓ����sW�s�G����N4�Jwi�@���ף��D �({l�t�WؓЖ]W�r��qj��p���ׇ�H�0�c:��c�q;u�MR�� V�Y/
)U�<�0��P���x�k�|:���K&m�<����7�<\���5�!Z������Z�~i�6����S��|B��X�d ��9���5�$�Ƿ�bZ�3�8J%j�`��<W�G�H�Y��s�/!s��뱄�Jm�{:�*Y�����"f����Z}]]߮"L�.`� �X�8�����)���Z}�d�����U�Ě��V׼(^�zp���\�PDZ�{�3n�dD�>OZ��eAyxs�X��z,���`�q3g��=L�C�3�@9����;��B�	�0�ݜ�<���R%�(.�O�01�&+ �+
(���zV�d��`,@�]r�~�ۼo��bS��UصP����p��\*�w��w���	7�/��h��u*�/���5t��E�3Y��T�ߜd�P�3��=��M>�9��ĸ.��6贸8����R��n�����Q��S���&�JsC���=P���DR]E&���r����lr�pGa2ƒqw�׹�le��JY����������Y����!R� ����2du4h��ٵh�n����q��3�b��e��7���N����$�ب׼ۊ��o�O��`���sR G���&�Q�H^���bh&�0��e�����bf_��&��bŭ�� �G6e�]7s�lV��&Ϝ8 �����]�N��.�G�]Q�g�N��d����v)�r|�C����4<9��,2��=�:�aS���!��r�)�?�����~�,�cJ�]�RE���Q��;�9�6����"��j����ٿ{4����Z��7�w�y��b[mGA�tO��g�}�T	��g����8s�~��7+{�����f�B������ʉ�*~OX�η��N�S��1	?�+��������^G��DP|����������w���D'k/!ϩ�g��1-$x|+���0s�Jh���A��ZЭ��dj�(�<բ��=O�����^-�f���Hq��o~^����`ȇ���^�)<y;�S�\���8�[�U���s(�r����O�u�*O�d+e�+ew�B�@�i=��2�Z,��Z	5m44��c��@��R�`��Ƅ\�3�Z���r۽Z�ﺁ�G�]E��C����2��;�
ޭM3��)|w?�JE l�8?l���iLiZ�l:�
>��7
>0@퐥E�Q����O+vi6R��\s�$V�7�����Ȟ�% & �\��]6;v�����t���R�^9����P$(d=q�?���&0 &#U����C��q��H��a�ɦ޼�XV �T�n�W]�pK*n	��	��Cg��'y8���ۑ2Q�g�+�	טd�b���;�JS�Y!���23B�2�!���ـ�?�AL�������2�X�X]�`�l��o�^*��Ĝ�w�$o�MQs�w�����M_@��>���!x���b�-����.�S�`�#�Dq\��+LK[{�
��� ��ώX�Ӂ��n�@J��	�wnZ_a�;ܮ���b\{��.>���:�X��ʟϼ��*�a��\��">}�p��'��|��9g�G�5E!�����3�J��[ȓqD00�vY|�z��5��3�oi��1� q���?�v~RY�h�L���x�
��,�`�tQ��"+� P����2�Z��{��F���O�՛
Q|���^���=(�w�79�����{�|Qx�ϼsᓹ	�T�lA����5��֢������lz=Ty�w)���:��?xp~��a�m��x]���@�yte�ت1>P<Ƽ�x�|���󀋣�C'���,Εh�i|�h��>"
�Ř;��쏓cG�X\4�S��.�0�&�)t���HK�tǽ

FB扎�,Y���f�{��/����_'����`��R�������}ׄ4q������Zʍ��e�|�
���K����mš� ���?� ���IpC�P�hg�J�B�`��zo�LV!�L��Pa��慻/�Tܨ�B�z�4y��=�G��J0A���3��i�`Ri��Q�v01℩������\;�d�0�.#1f޵�(@��� ta(����7��P#4�t7����1�4�[ߞ�`5�m�A޳,���+��#�҆���-Y�4��~kJ/Q�hi��	�i#ĐKR2ł�I`	������8�7{k�i��nm5������YNJ�o���:�[��=���]�-:�~�7k��^S��:�iĢ�Ŏ��ެy���S~��!�r�l�x��Biii����&>X��? i�"��UX��2-,�ܠ4�I��Bސ��0�Y��tQ�"��b��:B/�C�'���Ju�y�~���vA�����@:A�� t�h���4a�8+�Y�{{osk�뻲��Ad�o�H��!��.n�B5�/���v�|�t��I�[�M�o�+�{pC�+/��2ȍِ,*\ç1�ߣ5Iqi`_��%K�ޖւ�Qɀ`\sA,�V*W��q�_3H��EC8�S�ƛ�7#ڳ>��k͚���Q�r����m��7Z��Vs��9�a�<��xHtb(��&\�]~��^(=[��Ė{���[K��澍��'}r���,�~o} c2Ǫ�Z���9�L4��4pNB �u/i�PC��&!�*71J�8�:{��:hk��Gq-��j,}���h�B�e3;�=���V\��F�	[E>A( �u�}�d����P�,���J�.����Z� %��'�(⿺-bN_6a}��FnA�����k��n�]�;_��i�g��ݹ?�&g�ZCk�$��c�
�y����)�e��*tP�ZA��.��X�J��Ɵk�6ب���I`;}�߷�3zn$�Yv��6�%�d0�b�b�3w'�ԏa�<����*Y��]3ፂ>���nX����Ɵ��I��r���V���A,�	IK��U:@Z<�Q��Ut�A�5� '�T=�u����-��|+_J�2[��4$���n�P{�O]�1a�SYX.`��m87v(�p��	�8���5����K�Ѓu��k�e.��p�!0*���!n�A*t��J���g���jϚ>���Z��x��x��)�R�����$Q"W���j$!}��l�Ǡ�~.��f��y*s]�@�����T���bU��C��� #���<nH�O*[׺�5���-�l�p��k?�9��£A�4Q���?Z�M[������˗x� Zꋭo���Ǐ�����_\T�����>��H�<݈���7�m�  ?1�Wp�1��Ɠ���h��3��X�Q_�B}��eq;�u���b#�X��\~}
x�1u ��vQ�S?�2�*S�*��ܤ��5�%I�*J@чr���w]�uƧ����7r�O�ήO�Ď#g�
�lUur�WnlV�B�d�عfD���r�q�J��&X3�� CQC�6��[b`��A�a���\1ފ%m��94��V�߮R�s��G'A),��N�X�;I��-�B�yξ�"�faR�Q%����hJ�:o��\��%��մ���	���G$���_\ļ<���'4�et��ֈ\\�C|ܷ�@P⑕�|�ͪ�}_N��F�W�E�X� c��	^7�iGH ��Y�z-�)�*�K�މb��xds�QGǄj�0kD<�O8ޯ���O!�c�<N0k��|�	��J��z:�����J$�Z�m` �@2�{Ij��U���`�nh<��K������2��L��L����w�2l���Xu`�<)��=�y�"+�U���q�K@Z���I��âi�	�y�������KI���t�I�h���h�����\�6"���+2D�:�"�5k͵lő�\^�;Y����p�2"̍A&��2@h�G}����:HX9�������
�J�/s�1�A�q ��]9S%Ƙ�n 2�mZ񎙖�G����A<��E;��Ix����t��MВ�ס����g-��(����<CEK�B�S!p|��Iڨ�	���:븝z��4<)NJ5æ/���_��h&Ӿ��^RU��v�������|Gw��{&H�MN��I7������t��)��+~i{�G���X�R�R��|�����H��f��H��l{y9�L8h"�����&\�ڇ��������D��:88�����D����l8��R��ɠ���\>3��!�.�@W}2CB���؜���[Q����q}�N�1�9c@s?�h���^��j@��@����?ϭ��������j��yG����,���g6j��׼�߼��
{���Y���&�
���
+��ub�m��r�^MU�
b��ijN�gQ�L�����ٟ-!�$�[�T��t)�y`L�����"δ�Qp����-Py�h�Z����¨})�
�H�t�G���E�OLd?؛�M�=c�H�4l��6ID��5-B��!!������^k<��Ց���8���s��eL!�l0¤�{�P<ϥ���A,�U_'����yA�nB�u��o	p���0��.)ó��C�j5('�V����5���}�n�̐O��rT�Wh}���I�Z��r��]��\��j�K��i�f�i�ɓX!���]��faۧ)��uLV�G+��v~<��q��]��ff�]���hK��tź`��	��Q�}�ފD�����#��nb�ި��z���ҳ�2��:qC���2�	�[��� #�� ^=����R�@O�R���5��T����K�$	�x�I��GWC�}]�D��\F�pv���WS�jQ��Ј���1���<s�H����J���\%���~��]�"��
��뫔aqZSC?��U�v�ug��Y
��,}�Lj���������J��έc �s����l㬉��c*��HǢU�0c7y�YTq�+��ƆYw�q��?&�Vsc�.T>v��Q ˕n��4�F,qg;�'��55=]WN-����n4��m��1�U�P%�K����h8II�h�R`���݀*b�n��R�66�!��3���^s��ۘVz��ag��<	Y[�7T����=C�q$���p�r=A+�2,b�
̦����0�jrf�O�&TP�kmv��FI1#:�п2� #���Up#�0vX�A�M۷>��t�]�u�*�!��#j���L��5��si���7�1y��V.��a^��
*�c�����>��<E��ٲ���ԉ���>��;k�ʞm{$�4	h5��}�q��.������Wk���H��n��KM��&a��Ec�{O�#6]�Y������E�J5��Ҹ�8�rKmɓ
�$���}=��}��֗��;��\h�U���	�e�ڷ�X˴��^�~�@����t�x|~�����+����K1*܎UmO
Y�"hu3�ry���ܚ�={f��)xz%��ƥ$a���kU�afN��ds)�������q�3hP�[���	��yr��9%;B��.�b��Z��@�C����ux���T���RZۯ �gK�AN��1q��c,��F� _yrF}�7 ��C����:��܁x�o�'DQaĲ�	�xқNxEs��V/�����ޅy�vZ}֠�2�8��q�a�k�ٍЃ< Q�%Ĝ;�2;�o,Y��>�c͕��\�~U�}�.q��k�[�2���~bb�N�����P���e�2�W�}��"��qG��>w�n��1�~��L��������(<z���9������()m%�"=��nhTk?�>�%19����>��1��bI�&��Htm�hp=��l*�����w\4���� "��Kˈ�� �8}��{�ZjÐ�1@����)� m��.�	�"�.��\�E�\�#�Y6<s:<��C�Ν����^iX8T'C4����V���$lOV��"O8W��߁���m�{Fu��sc�ƿBXˤD-���t��׺>���֌����Oi�����&x"��!��qk�r
ꯚ�q�9Z/�*���A�|��?m�\J��}�"[''.!�����옒�իUUB�4��,	�y�YL�e�:��C�=���Q��ӵU�ׯ�(�&,ڕ�'zE�3���Bq��mH
����[W����+�1���ɕ�w?����$�@�����Y�^�d'��5�������:ACj�5,�q���n�G��Y�u3_��)����N�����ݽ.�0����!�If���1A�,x]B���p�A��P�[��@�ļ��~({z�HC���m]]�O���u�p�i�<�u��ѹ
�%�P[��ei�A�@�F���Sˋoߛ.�?�b~�5�p_b���UU�:UU�9N��a>��/U3�tE���;�U^���^p�����Z�wxu�������&�t������h�1�``lL���Z����t��u��|�a��9�c'�t��d*}�,�G���-z�<xWd}һF�5�˭����T��gO��E�#|����ެs��\�&��K��O��vzR�9 �<�X��w�|O
��z����]mf��԰;�}�X��	?��x����S���B{����7�S�hy���<2��ҒKe�nߠ����,�Rz�M��c"�'������JW勮�%���b��z�g��55��8�؁���an��O�$\f���~����ŭ�U��0�fk*��%������N9�"XK"�Hq�DWD[m��=�S5<�y������a4���w��޿n�vr=j'��t26;��ך;>oڌ|�|���AL�R�&������4,���ԄgF��͖�������3�+.�G�=��=E�RJ{ٳ���h� L(�${��"�����͓�*�f�x�\�'��u<*.���p����s�R����^�㗯��s��.6y"�+
=��˒!i=\hv���ULo�Qq�"'pl�����4brS���1�}˭�RF��q��`U�9vԩY�d������W�?��U6�s�'�4vvw1f�����'���y�t�.B�O���P���^(S��փ�Z>	S�Xq}��ڭ���a�AH�%C�[<��.�G�N3��\��,�X�Oϐ�O���FEJ�A�M����L�:eA�MM���&�#h�h`zB��Y�nF?YrN��\�*|8B�+U��9�k�c��[��rk�o�o�r�1I.�S$S3�`�:��)�W���w�6��'�X����pc�+1A��k�,��,*�1#|���m�>�9�����h��nB\]���bM�'�ݠH,���}��ِ ��`�9���\3*�p��jB[�	��!/]���E�ȟ:@� �	��c��z�+��+7���t���o�"}~��7t�h�y����&�������H��æ�k��F�#��pm�I(���n�mK�A/���6��^�1��{��Y��w�m�h������X�E���M��<�����s�痝���,��#k���I̱��埥���h`��1�A�ӯp͜H�����������޷\� ��A�P�X�G��ys�������^t���V�9��鱯�P�2u�d32��?��r�^/��,p�sA�Q�[�c4v.ʞQ2�]'�t��fr���y��Y�l�Ж���J���ql�RQ}�mէ���bM
�5Y	1ɱ�^��!H���"�Q��rO�I.?f���;ܕ���Q���n��B*�^���Q?�wT��Ȑ�<ĵh��znd?g��g��v�ˬ~���U����nm��Ы=��v_�`VD��sW �c�����7.��P�7]���_��zX�
O&o_��QW?��.������ꠉ�E���4'_���)�E*��!��X(�U`|I
��b�Eˆ<0O�GY���?HG�!�V�l�K�x��$�~�>��"ӳ�����
2���e���&b5������C��NvA�{������c�Q'����G .ڝ%_���Z�K
 *��I�Uɦ�0��2ɔ`��@�"bq�Sd����5��6#�`�(�����C��]::ar�T��L�}�JxX�G3{�᲍|w��#M'ړ�i�;"ϝ�� ���'��S���5DP���pj�S��<��M���ǢY�(�'�e�;N1��l9��^��m�C�%A٥���������R����V3ˆ+m���mu���<�GlU6\/7:U	?�0N1���������[iqy���X-���Ǐ��r�`KE���v΀�Ix���9Ud�UA��z��*M�g�o[�oL��&v�9^hL���,�n�*�}�:_0���"��|k|�˴7r��ik���>Vc)�hk��b�G����A�b��jP?�\���<�H��7���^F�{���}��`����mapVm�e��Ɖ�д�%�aVs����_�p��ݷнm-ҡβ�s����H��Ӽ��_v���t�����"�o�M}��a�ō$ѱ��f��n ����9��&+=�g���ղm��PI:	ƴ���K>��I��3�慻�rOv�@����t��0<�|J櫆�_F웾�5�#�!�t����g6[�f�Ҟ�#={�]-�G���
 ��pX�9�X囲�2��~r���>���wԑ9Ӫ��m��l��	q��,��Z�d{�\t��~�;�\J��9#Î�L���f&\$�{ʢUy�]<�@/��n��?4���j��4�����j9S�^jU~�t-�' ���Z��ݡ���l�H�8_p�RZs�>�L��!��CG�
�G����_5��O(m�**�,��Nk��'��hp[�����í�A�q:�B�����\�g��1 ��k�o����Z����Q6����(�Ŕ( � ������5X<�Y�ݰ�}w�B@v3�X|�G#|�9�>Y�q����x̲��;��ݽ*�~W-~v�q]b�ݻ�L�)�hE@ת,QP}_���/���X�'�u�<��t�kP^尖�'c�s��p�v����.�+�v�m��s�k�Q����!�?� I���则3�u��C�z?��fHRb"�oߎ��"o#ھˆN�	s��yr�<��ͦ�����~��{�(�pRdzS���N�}-K�^|��^������B��;?�O>�8��S��U������YR����y���myE�]��G���M�HA^�?��Q��I4Gq��{T�5F9� �����c��-c`Th�[�/.&�����uMc�o���͊�R*��QJ��X���Dx�oE����mZ,�2����'U؈���,�1��q�5�`�#P���n�;jTq���Ȳ�Ĕ�n�]8���j�<��7EE��y(�$��E㼈5.:.|�S�M�1������#��f���[�S�� ���ϕ?�Y������R�j����R����z��gq0#B'�y6���N<��]i�O#x�N��9��gԴ_��@P~�&�3��%�|�Ҕ��������??�F������ə��LEl���ׯ_gk�Y���`/�|Cy�l�ϟ/��ҋ<5}&�cyY�E�����Pz�eDS49�׶�����A�j|�5��f�ú]:::�ƅQ��)))�53��ƳG3��?�%�3�K��Dwww���1�'�ݜ�w����R��i�X(sM���e���|���Do�R%�*�� �_��
���acZ�7�������lS(����d���w3-./��L{����ף�v�m����89���G~~��k�"F�z$�h��DTTd�
�ڟ�}����@h�6���*�=�#ԭ�9v�i�����i��1t���5y�K!��5�����:'���O���|�u�up8<\I�؜��VO��ko^�lK��m����ʢ���ĢJ�V���9���Lp)-ՙ��X�z��H⊢=��4V����֔��"�$R`%rww�ߍ��V&K�k�B�Rg�Tq�׍����&c������SyC���H�O��R7Z6	޲��x�s�z)�PȲ,,-uM~�"}N(5�����Q*=�Q2�Y��u��Y[;|��#:�\\6�-�*�g�����w9p���0�����
��n�@����8{���ޞ�	�A�3���5�ʏ�Y\����̄Sv�L�n��s�Z���<ecc�&�r՘/4��
A�����o��q��HEU �� �.��@�=m��STDd,�4�l1[)��ɀ3^}�������!��֞��l�y��ɩ^��^��G�d�?N���%I�
I� �h^��-t��k�G*VyDA��ƳR����S�ܸ�����j��b�Gѭ�����[6/<jݸ������'�4��eI�{{m���u���>�q?��~����v��7+�~��3j���ڪ�+/�&LM���xu8��2�("��sg[�*�)^ v���Dh PR���mұ��{>i7�������C��8��8;[�])P ]�+�>�\s��q�%	]�`iD�D
��Tq�~rW(b�j�P�a��X����F̄:銌��I�"�u���V:4%��3�xd3~D���xA��ȤB���&F�{Y�r,S��޻���� L��6"�1]���aE�Rb��A��� �%C��`�#%��>��I%��^��P'
�11�y4SXAWIkL2-
�$�#r_Z�t���X�M�����zx���@^�H�|�%ݮw�Y��m�} t[f>�+�d���|K��˧�����ZC��pf>n � -Y�
����I$��c�f�7u��uZFQ�2�h�H{]*�ϯ|N��x�ʲ|����_�]J:�#+1?�f�����^�\HZLO���]�x�|K���� O��"�l����}���1�Uo���J�������o����������I��o��{�D7}/�`5���Hr���d�]�9HoE�q��O%T�OC���ꅄ�:K��	OC�f�7� _S "�������ӀY����ub�D����LEF�������׈�V�a2�����ΰ	C�������}�I���p��+�A*���ԘR[�.��pQU���|^��e�E_���a|�I֘����P�[�~�4��Ĝ�G�X�>[au5R�9�"�bsJ]�B�v��i����¾��I�Uu�j�
Q1���h���������r|3=~�Y69n����8�B��Ԫ�8�Ņ���۹	Zu��|�2mjTnZʥ��ɳ��&%B�o�[��Cx�p[|��p?�������m�m�]����QНGF�A��b��w��{_��)�v�)83���2�ǥR��n��\������e��X �:=��x˄Ý�"���l��xr�s)�GF����{{�Z�.�ת2�Gx@�N®3�|�a���0����͝�g_�;�B8�0��o����m��Ǆ�$KZʐeT���R}�5d}1@�]8<�uF����߃:B�(�Q4�9����,����?�[��H�<��/D��3�
n2A����J�LM}Ml}�ܷ3�sr
bŁL��~�9e�\�+��o�LX�&�6:ܜw������8âv�䲵����N��'���7�q"^�X5�1����3���Bgܘ!�:�av>�,���7N���B�)�@ѥK1�\o����@�N_]aݔBh_C�v/7o�y�k�sz��?O!�.�Z�;B	���=��&Ukm����ynC���&f�� ��~~~=����l�����*���[���I���=G��P���%�7�巸?W~:Z�>1���� ��l�T�k�p�ت{�Dt�J��[�'6�jC���w��1c"\�@Єu*{�&�]���*n)#�)q�}�ɼ�~��ʲ��K趏��9d>���m�]ʹ���Nb�(A<���7}ik��^"�Xș���J����A*?`��BvUV���򗇼NuY��%q���ˀ��ӫt%B�H�y�J���@���Ⱄ���?B�C��7t_f�kS0��}�z�����e������%��JW0�����E�u���������:d��9g��6
�)͑��icŀĂâ�Db�����N�5��Ah��ÇKicc�׫B�?c�"��Oչ�d�E�C;�(>w�s�� ���u������u0�<c$�SS@�D
 &"T���X�sO�M��Q��ב��&�[�(Eߘ��.S�7���ӷ2��[5:�9��������������9s�sgӺ|	5�Qb<Ak����nh��pw&������~��V8�ҳ��r${�w^�:b�����p9(���#�A���9�5a��0�i�W}:��cx�݈�72L����o�B�3 �ά-1xt�_ۦ�Yo�m����#	�ʖ��G��.�F� ����]��\�4�7��ׁa�aIT��Y�z�|r��jk<�}(�22�����F*��;�}}铯2=35i��V��?Xs���@��Y�t�����'Jh�l09�/�Z���o��_��� �%��AN���Y���^������2��2LܠK =� �O��lV�P�L�����_���ʔ�-���%��U�\g��?��Kv��-�Ƽ��EXc�b�̔O����f�h$
��Vjp4�2uh50BǢ  1��4H5�}��`�D�TE!�N&��X��l��o&�O�F~����= U��AC�����J�~c;�}��
�=�y�>�2�wǲӀ�Z_�]Dr(M�.Y��u#�2���'�R�y��<��OQ!>�Շ��M7o�3�����������+B�Dmh5Zm:8����X�����p�跙Dn-�:��?�?O��[��<ܝ��vFHt�����5��hZ�Y�R�'=�溚ۭ��p| ���Yȫv��4~
�ۧ8!�x��RH�Ăv��g?�.1�sF�	N�X����.���Dn���C,6њ��|��ֳ�.���G��e=�h���oY�m|Hܾ2�ު�%���ݿ�&�V��V��Y�{A�srq��lh�E��1
rY/(��3�56W��I���ExL�;\�H�Hbbb��O�}i���?rPg�`�݆���U³Bi~���pI%%��]���<����32E����V�R�7
�|Kc�J������k�Q�Hh<D@,��o�B�/>"��V�^e3o���o�HSjo��<|������2ڻ}*lĒ�����1��r��hh���*����v\ r8O}~ܨy����S�MXb�k�����_��/_v�c*��~�:
q¹���(~��|���ϯ�~����;a�ML� ۓ�j�aT1��W�2����9�Iѥ\~_]]�Ъ�F�L��YdC�Z���_�ct�g�,N�����Q@/�nj� m�6�qP@9�HFEF�t��Z]ݸi�3��w�$���ŔG��Q>>�( ����I�+ub��锫��]:w���� �	/)k��%�U6yŚ�-�4�M�n�B.���6(z:����9���n����U�#Ifu�>Q���v?�Vz,bTN�r�?��2*���"�%�-��)�ҝ��)   - !(=t���"���9��s-���9��}��8]U�������8Z�N=��#X�u�޲��ku�e�/s�Q��'e%|��c���C��2���h�YP������J��%KʠU��C��JiP��:3��_�yu't��� ~���X�>9�V0���z�h����oT��Du܁��^���{�y̔����1t"�jҎ>���-O��\��ѧA���2,��]�w�ص���I��á3��@������u��M7m���״2�j���b���ʼ����	�����{_���XI������JWy,�Qa�}�caT7�:��H+�.ueM�#�y`��F~�i@m�a��ɐ��0��zߡ@.z�Nf��VҔ4Q�u�Y{�y�rQ5g[?5��t73���K.�m�gY�uC/|IG������,���L�?<�-9$hQR�����c���.���%�������מ(tɴzƩ�"p֤^��Ӡ"5��C�]�D��!O$��NVI��ǻ�M
#�lz5�k7�ji-}_Ry��/4���C'-y|э�ᵈ�2��dnY6� ]b�wh�rJ�9^	���̈H���!s��7RCx&U4���8X㕚L�<�b#Y�<n�5-T��K̴h���vƩ6�M��sA��E6>7�Ȳ��g!�\́n�_b@Q�:�l�H8j�ˮ&ʡ��>�W��c�xa.��jj����{ �a�N�+�4�Mu~���Tm�/JM-:L��M�[Z��O��Q*�Sb-���/0���R#��m���4d�&���oBt$�P��n�~���'�=;���E�ak���]Ր�OJK�_F��s.�C"�-?dg�ǯW5&��-ׁ�R�� K�}e	����rW�~u �p��(;y��Z�߮N�t�2����1����i&-�v���z���7U3\)�sy��L*ް�i�4��'x:>	'�d8=����Z�|}��17��#��+$���],�`�㗃�ߠ,��� _��#{����ʓ?��z8`^,YWO�z�������׳D�f|������(�ZW;:���f�	l���j��dy|iW{���T��ѕ@�a6�[~zb��?��9\T��\4�ڵ�0j��nb�hH0���b�C���ĭ%�����k�ј����jl���°#��48����uAK5J��b�cY4{;������ikн ���U�?<�t	��(��&���4"v�h�
�^Z��/��ɣd�>{�tӃ
meR�6�4��fԊf.�]��%@��m��4��3u%�L��x�o�{������d�*���r���SY��iA�0Vpє+�Ww|�ڽ��z-���<0�/�E�'����(���`��@��"r�Yؘ�,֠����"Sr$P�s����krK���Qy��!�.����8���b�nq8S@�"����g��]yS	�t).���{��_ʜ����-x+�v��b��n�X�4�W�8 �����>�*`�n!�af2(���1(f��
P��]�0+&�m�I�n4�d�b��C���.Կ��,�����*T��~�:�7�\�Э��/_�r�r7����;����o�h>���I�����������9�r;�O'�?	�`֫���7��'f��c%Q��Jb�:��U*p���5&�<��Q0(##τE�h��,�h'3�>S���˗/7.BCA(c�[�vv~�^����r;���������)�h�=�8�lj�4���9���xY���糝�l�r�|�AU���_�<������ ���־(D���K� ��P�bqwPO�y�{8�k(�i5�`*�.D�299��"ZO̍�[�Y��B�sG�Q�#�0�K;�|�5�:�=F���L--�WuA���[H�Ĉ�i[7��1=�{�o٣��r��A���Ɣ��X��������$2�$�z\$�I��qr����Av��w2H=>H>H�(��:8��tt��a0%�kiq���Q%��Bmb)J�Gu���ڬ)��R>�����2s[�@��Ah%�ڐ��X4�S��m��y8��}�r����'Ko�M'�a� �Q)#.�̿�8d��G�yv�Y�x�5���GQ��y�[-hV_2F;!Ǒv����r}݀*55?�Ś6E=V+r�*�[G$�L(ߑS��)�i�Db�~"�)���."_���܎������0��,11���� :�!�����-�b��W[[S��?Q̆tr��Գؗ8�E���<�O��?Z��~}�jV��)F� ~��I�;�U�+-��(U=sr�V�{Rg���R�V"�hd~�֬��Y?�S&�Y�绣vX��F�����ߙ�"#@��X��8�Б⍛5q	����a��n�
KPåM��R��K-�iݜ����F\6��������>.Ů��v���BFYb������4� �H�$B��A�d�� ���=����G����)�3?��@w:|�&�̨�q~�Ov�~qOnn�	3~�󊿂,�t�)WK��=t���u��*"�6|��^:R���j�k��SOӝ���A���2�@��p�?c�#�_��c��H��d�х�b�x%��ʝ6H5J$J�-��D�z��BK�;�!���� gݭ1~��ʑ��@������,
�nܰ�Xl}|������e�%�k'\���4�����|L~vW��y�=��<9�E\PS�EHq��G��ÆooXgN�r�ܸI�) b�|d�2�kF���|:��Wln�c����_A)J�͆�Fz9i�"dZ�<���G�A��3�r1D�RX�Rʩ 36vd�c�p$�U�u�j���mJ��-����.n<	`�����XoDozma���~K}{�!	f�O��d����.�0%�#I]Y�T.&x����yA�����C�{_v��NmFaٻMuאw�@�?�$��l�A%��)ה�,�7k�t8M��"������&毶������4��ڱ&6q>K4·<�jE�Z���בp�f
X����a�P\s��� ��B"�Y~���h���"�k>�^�']���J")>�i�&��Gh�?�i�^��5��>���-�O_��t �]�t��O�f���K�I�"�E���#|����VO�6g�L�P� IG^�_���kg�R���4�V�r��#���ۃ�F̘�|�Omՙ�k�k	��A��[�����pڏ2�o�:'36��ZK;�5 ʩ8��2�WL�8q��!�a�UK���P/cGW9�1=A?X�	l�+�0�n���ļ�(��/�^�5#��'��n�H.�'i �m���I7�7��fO�>wX�<�Kd�?�w����/(���[���/	Ǽ�ב�K$���s�����G�)��K����FGGG���u��@�[)�^>ջ��2�D��������qv���J������Q�cdJ�O��M | �0To�f���~4�mv�-���o��Z��N/|D�l�s�iH���%8Y�س�.�:��\`�������p-�Nk>2A�[$SbC$˼l�-�ml�R�[o��W�K�U�C��\-���]V��V����������H��) ��^����Z*_�<���'3��4ߑQP�Q#�����d��e5Z�xB�w<�AD"�:9����k`=qs�#s�к��|�\�b�o8`���,E���[�Ja:��~��N*vB]
R����(I���ɩ�⁪y�q�*�.�o$=X�7Ro偯��-sx3�V�vҷ-v"e�/����^�LT}�B�JOE�MT:$H�1f#j�A���Ч��Q���W}��� �>���]7�S�e!U�T0��O�4S0�Z:�sd��'�@���^�?]��%�O3����cL�f�l�'���QV�r��&�Ef��Ԗ��g�t�9�q��n��3��8�&+���pEq<{]�h"0�8�1��i�9��tK��!���7�5����effV��ߌ���4����Le�&F�=�nklL�rN�����9���:�}9;>��]t��#�p{��Ȱá�*��
�E�|� ��J���M;����k���ڸ�)�`�z�u��UU�.z?1c�]�(t}�5Xr����pc��6��>~�H��	�_D$AL���wM��{e����q��B5�}lʄH�s�æ�+>b�U����w�+�xuK�J�ȥ���m��^WW�V���K�;�oØ)m���U�����*��Q6��2�P `D$�
4%�fDșO_�ELs��Or�X�@���Ei��H˕D�����O�E�(o��:F�C1]���W�η<�I>lJL���Y"�[�x9�{GGoO��+qv87������p�s�6�� �%G�k�pJ
�px�������<���S�y�k������Y���ԥQr�yI��]+j͚P���T�T��*;é��(���R�>��S��]K7A�5bg�GW���`{���46���J�����!$~晘��C^�X��a�D(~��)ic�)��ٳ0�����j�'+e�3j9�]NI<����x:/l��i�\]�v}��O��<;;� so�<\L�-Ķ��3)j�-�?�?�g���4����XSP���~J܈5E[Z��M�q�w����t�4�{A�K�a���?����]��K�-#*$�R���^��v�9,��9����
���i;�����8U��� �5��,5��9ݻ�Y{�o���������/�Lma�����ʪ���V��	��vY�D���_�|twQ��z�L�F�?xDP�Ӛ�"DV��̉�ԥu���'+�F�8����%�t~�i�Ȋ����N~1^�l����`�7p�C4]8�	�AB9��\�潆���+
�9���(|�_"���W@Id}
M��>������kU|XP#�񌀮EA��@�jU:��I�E⮵
���1�^ab��] �466�.,f��e��1=Ɂ^%Z����/�H|�!�e�K�h>���!����ғ���D!�a��C��p�%O�n	֬:�C�"�e/^�������F4�1������"-V��w4���8d�������_6�`l�A
b��j��zf���g�g�%3�ZS��I�<;*L��(a���C�%�`�q���ѫ���׫��/Tb��h�l��W�m�t��0cp���$}�䭹���'!!O�Fh��,�B��;ߒ�_�[�w=Ǐ��2~s���g}O�pc�H
?dT&��� |#����lǀ��%�T4�����kp^��*���^P�5��t�@��t�m�U��_��8s#�V����D1g���{�kr�1�'�o{x|:Cy�@�|�wD�����ѿ�p+Z�9�I�`&��w������
��[���O�}t�Α���F�Y���X\�XjQ��뱞�F�R����4��-��y�~�tc�1��-��#��'	[^���<����������͙|U��o>.�( ��6|d�>;��ۦƸz��u�e
�bM%x���FFF���5� �2H���!>q�V�WG��@0�3S���NrA�VC֔�H�7��H�蘟T���*Z�"�g@����� ����G ��zU!%Y�&W�QX�Rx��=��_5	�t	{�	��0�E�`���K�{���p4�gT���)�>i�5��{�K���U��U�/��B19��-�K�đ3ȥ����:eh��7��W(��s���wk%7G��)�>3�<P�-���\���-_�A���^���pc0�e�?P^],s��˺�1>�ý�[�D!|6���>��o�kAD=uu�([\��G� Q�k<�5�l�-���?r�,�P�P�p�e� \�ʸŷ��`�}�M �ݿw���0Lq1��N*.f�3.˓�}�� C���ڃ	��<����#Q1�:�v'�=�2Lӵ��KM�����r���~u�̪����-���wSc�`\q�N��w��l�lB��zq���b��г#O�t*2���'A;VI����7��P31A�����Ce�V��T��-�~�~��g����eP&�бvv欷$RӲt������%�H�z��x�� J�,����Z@�J�,J��K��CTjA���Z�aUwb�m��Q�(!����]|ݚ'��L@i�%18f;�>Q �8l�g_�><l�$r$��-ƷN�:R��� /ooo����R�p�*K�A��~ˆ��|F�T#qw�'Wy�>���.V�\9���B���K�����,����M�*~)Q�H��0���P��ol@����ź8�-�}yq1LFJ�k
�e�����^�e�ň�U�<̞��r�A���ں�*�*��ጉ��{����y��Ly�S�uTİ�M�{�	�%I�cم���-��(}��>�ǾF���JQ���dL�cP6J��
Wa��: �>���;/F��@�?B��v��^�r�~ &�bud����ր��4]��J�7���%
�����>�k,n�="�:��=�Bs�V�x�^��f���_���ʖ)��R��U�ktA[Gw�8����5C�W�u���(Kq�k�`�i#��HxvrR���v�����-v���WDD�P�y���j"f�&����D���j0�޽q�2\��͉Sc�wx�"��	}��,�)����m�vt�4c��LKy�̙j]6��bn< ���iX�f��Ԝ�Vf�>��5���U�Ya���U����o�0�,N&eh@d��{���t���M��Ae�N�=��u�� �!{K�Y؟#���&��W2w|!��	�JG�M�[�&xЪ�T��]�����犇�v'��r�}�L�8����G�x�)�B��1�;Q>���}$�l�.��2+��o�p��d���w��r�B!��W1���sj�,�n�Y��r���t�6}�w neB�L+Z�\���r���7;g0����I�|�zDx/ڰ�Vq
������R����T�m=?D�:��c����XC��ڨ]�C{M��ȼڮ	(��$��ޛ������?���?,=�}.�Һ(�w�����.a�Z�]LL�B6̷��$J���%�S�=Y�9��UY�A�s�;>�O�l&����� b�YU�䟹Ϧ�pc�o�a������]��e�����Y���/�9�>�s�QHM=%� Ғ�[ہ������?�n�^S��� Ρ %��ўXfG+aOLs�~&q�3_2�Vp�_Q�ڵu�\\;q��s\i�����vQ�Cԉ)��o�"�a-����J���'-ˑR��确���'w���̹H�8Ҫ�Gi�翈B� p�b'<��Ѭ@G��N�;�� lV.��,�L��П�_W_�T���ji�Ѥt�r�Dwt�i�-PD��^;��p���}^%���߸6TRGg*������?��o4�|�w�4�&�B�5q@��� _�olC>w���!�h�u[�L�e��l��q�Yc
��3��u?����<�CKQ`h(dR�^]v�ZH1��W���H̔�8�c)����r�III�S;wp�����b�[�c;�H�h��ձC�0 �w ����s�z� -�ޟ�g]g�E�8\f�V�0%:���t�?��*&&fz�Ӻ�HT&����e����z��t�8�֝�xL�˷R�^�:?4<<,�6GJy��`/�GJU���V�@�ש0�=G<��ǻ��I/��q�(�E7c]qY{�M��o��u�:雉^��љ�D��C�n���@���8���ϵ|���/sp����[#�r*�Eя;;����D��(K��J�,��V>}|�B�|TF���v��|��ĔCj��`F�]�l��ӭC�a�?��c�C�>fP'��Iv�eƗr&"A�
 NA�6|AZ�mϽb�����u��\�b�V�t,�� ���E�A��͞�xB{�!�_��;~��9J��<���D���	��#�-�3�u��<�/d�#J����HJNC-�c	~�4��P��@��0F��2H/��]#5k=`��53p��!���-s�#�y�;$�'��7��T�g��t�}[��G�}:�W�\$��/��Ջܔ^��F��M;�w��@
n�5��O�~�}ǈj-��Y5w�3妵J1W�cHy|����(�$����Tg�p��6�t*��m�H1�t�s	D����(Ƶѐ�X����B~lg��O�B�cc_�N�`��Q>�F�{(��ս�Ǧ���kc��]D��˥�Ռऄ�-����Y\���B_K.�F�2�ě��f\7��R��[��Ŧ��/*��)˯�ܵ��bO�?lw��0e�_;�}�qX,��tq9�}�z�7?}�1.έ��x逑&ﵚ�g����C.��`��i�G�N�Thi�=�3
� �����Q�'K���:q����iD~���I�<k����)C�>\ ��4Aw�|�[
p�M�x0a�iԷJ���پ~=ι��-L�Z�Ö2`���bji���cT*Ǡ���K����gM�e�VT�OLLlF��	�
_mGW.-�h^ �b��ۜ�0���#{���<U4œ���a�>����G�F�w��+��3!�E�C廂q[B�+x��m�c[	j��-������&C�\׻f�ߎd�og^�;eg���1
H��nɕm�����[�W?�n����W�ߑX3��f'�`p#���!�B��JE��"����H��K#U�Iصr�	�/�}��d8FSѨʲ�;���=��y�%h41����R)m���w����Xz������n�!@��xyz��F�)�;H}�j�?���5������}�k��1�Y�k�TrK�6>�t�m���h�Q������Mާ`:�(�����t�'FFF��lj���a��f�}��66��Uc/�7����}Q��*��:Y��(U��ٍ�bѸ��3Y�����vb �������r_��W�.AvUj.�3>rȥ��1����@pCĤ�!Έ|���@a?U��(Z6��n;e
�.ϛ�~�{�쭘>�ɹ9���#	��_�0Oz77'��D溺�_<��\(�Z�c��=�#~����M�w�qaI�_��zfQ���8���	��yt{�{FM�b�Ư(����%.�m�[n���D �b��"�=lM Ox./,,<��-I��=Yf@]?�0|��d,U��p^3UVޭ]�SVXR4����T`��U�Y�^�2�DN�P��?�N�p�3 ^a��c��Ų#�x|D,��J�F��Wh����+5�����������$�	��r�$...d�t^dc<��kj�\Pz��]J�_�����]�"����ֳ���[.�F��
��&���� X��*4�h���h%���$Yw�8c9wwB8�B��M]:]'
Z����lLxY�I���f��6�}�仴44r��u��Z�E|ڌ��1B0��%�J�ׇk�aIn�E1��\���	����s-�GF�:	kD�ƥ1M�i�":"�9g�6�����V��҇=ޯ�>ά�Ԭ=�H��M�h���I8V3ƃ��=��߿k�%D�rG6fk�%F��ϐ�et���!��峛�ۻ�`�����D�	Qy>��W�q&Z�Ǻ mX@��{��JOZd33�Ϫ&%&�N�[�5rs�!k�)�k^���!'2B�7-�m�cI�1��[Y����>荃@I^uZ��p��q>{�x5��i�^�Ω��������y���:S0n�&��V�`��輖.�zXCF�M6�W���fG�����y,�}�e��[��`�}� �8�z���www����bA�.tڀTX�(�.�Ux�v+`�Ǉ;j�M/�0L�˞��������Ņ�KV���1�&VH��U�ｋ���I�_K�Kڊ�omK&�i�A�����g~��������b@��3(�{M�؀E����InR ǂ�$�f�-����\?+m`G�G��qw<8�f��B��kN��lT�[��<�x��"�G
��+���,��f���#~�����F�^Ͱ9s��.Vdڈ=f���}��ҷ�]���=�8TB��t���b=v�o�S˴���K����H O#�77��^(E�L��ss|d�mE�����z��؉�([W�hY���DC�ifn.�X_{A�E�����x�����W#�����ES; ���$T�l�]kL�7����ox�ڗ3 o��g
1�K��c�W��h|�����QgCN�оȈe◥�QT�]\��,����N��Y��+�-�^S��"a���.f�|���<g*���H�ݧ~��s�R�w�wb�^��oX[��0q�|R�mj�M�3��F�6�q��/�r�"e*,�1�1��R;V\-��%�E�_�	��O��'*��݃7���v���E�ŉ�/1�=U�����`]�^����s۞�'/�p�{]�&���&S{�?��
Q�����Q
��A0#���a�U�(O�k��Q�~١������O*�hܑ�&��)�Tj��^�>[���u���$����2���!XK���ew�X# ��e�H�B^�\3�������h���3Ȃ�6����/�=�ט���f�\��ϟ�`����������!'oQ����ׄ��M�;T�����a�	J�
�!��jP4��U$\����g���of*+�_ǣ<z��
�'�i���}�D,4����^�k��	\������_W��V�;m/�;�Tmhgo2���{<<!��Q1*��M�"6����a(�������3�)�a���\u�ν�Я���:�'��2��/�������+�u����ć��{E���(8T��K�[7��Z�2�Iuxn��+�"�[�6}֙ȩ�z{�G닯�'J��C���^=S��n��x����%?�Vv����QYa����#Jrr��	�����VU�����&�,��Ŷ1u��1 �('��.}[$��<{��N7�D�9P�;����_�ЮC<2L���޼�ռ��i A�K*���G�L��}� >mY;�q5$�2� C+���`Pl2I�6G�-�mC)�E��Ө�ro�3�hY[���C=��{��7����& ��g!
q1RuQ\��&�,�+F�iP��q�T�	���l�1 ���mf��{k���N��\\eF͛�_�S���~c��Q��ñ_�1T�j`+[�WQS[Z�S�����m]�
h��Z�g�ށtɊK}g ]&=��W� b���w���L��݆�:Z���t����(s�a2:F���Wr���^p���sb~A�">�d�pѦ�,���˔י�Z��7?�X�s���<5B[(0���jd!¿Ņw[�=<��"�5�p��`),�Ge?~�0T���n�>:�tk4�D��VH�~��M���[N��oF3ᇓ���0>��㬚�%)����f���,�.�QA�_�x��uy/IX0�����rT�ux���bo2�c�)�$����aC8�,B*�ۣ���0ыo�><�C}_۽���t���.�|Dq��T�F2U�P	����g������B�n��/Eh � pK��V�dXK�_':0U�Z_�5��Ǔ����Μ]g`�7x�D?�'&����;��a݅��SRnD���n�<�X]Rb��{+��g�1D� Pe�ayT3o�9���{F���D�%��^K���񝀆�Ǹ��B�@�t��Q�	�q�7�	��5������䅳�"Ñ�/�٭����`�!�a�R������$�/���;��=��G4�P�:������;8xڃ�ݩ�������)��N� #�e��{�!���Ӆ�/�-F�rb��zV� D��DEE� A��]wpp z�ʵ��ۘN1��D��0@_���b��E�T��~J#��PM�[)�6��E��״�q�D�?��l��!�-L�>Q
{��'�=����?���J���}���WRsp��2�g@�T�x1��y,~Vzm=v���[7�c^�|�cc��V��8�=��̊�픸��'&&mF�dM {���z�:�c�{j�����X�F���M�>���ʞ��7g��ol�������X~t2*���C�\�>�o�k��S��w��W��.�'u nn!�Cpt�`���V@vn���/)��u�T�}���o�0�!�E��c4L�n~��$;U�^l�87$
������l1*JJ����9��2W0���b[���./ev|����4���*k�Xj'�}���a��(���'�������3Bd%��<�FFO�|˓�`����XPf��vv��{�ìJ��\g���~��Uچ5��������XTX������/��F2��k��,�M��o�o�_ӧ[{��gҠ�~��A���'ؑ]ೝ/&Q��Z��3�>���Ғ��Z���6���\R�?��y�, Lg��xY:g��aVkq:'�I���Q̆��F��Y����a�T�¡�3�p��upnXʐuu ĩ>8a�8:��1.]��u	���2�V�*~�"D8=ġ�:|>&o�45YnT�~V�:�2�G�.�m����Nf>}�hj!���i�ag�"�dIB�����{d|Ҿ��{<r����B�M�u�m�&uC�A`N��������0�i[�IC��du!���W��m���k�:�S8��޾�>��Hdqxb�����}��ѯw�f=�/.jA}�c��Kt�0u�_�|y���Zc1p� -;b��W�p��O�P��~��5.~�p-��3�R��W&&��-{��᳀���������f�.�/��(6�-��`�_�3��L�D�!���?lk�����AA���h��D��=1v�x��Re�(�sO���7��hW?x���BI�ȮA<�ّ��`b�8҆q_U&t�����.a�e����[@.���D�Z]��"[�=}�.���Z���.YDk��t���n�\G���L�O)���n����`e��s9N{6��sMU��]�^��%��E*���R{��@f�< L�j"5�#���@��v z�z��K���9��D����(���dBW�$�hܗz�o��O�����s�uؒ��\[`h�T�ؤ���I"@<X�����-oLu�+�n�Ň��(�GtD줛`>u83ߠ��z�2ޅ�S�c�B��R�g9=��+Q\�H5�����sQ>����;�kNy�:>�˂<@�T��:��O�A'l�x�k
>�M귴ww�Φ{�B����ϯ^R��:aX��spe�%�d��3㣵t�<j����?!l�&�g�Y&��-FU�'N�l�5����pŸ����L�\���O��a�6I�e�jK&����t�.�
�1��Gm��'T��r�/.�J	&'#k�>�
�Id�����-��T=#�kt�%
8�_v~�
;.C��XH�m��q��7ޙ�\�����券,�3N;�z۾��H阓�0F��qv�E���F�����ΡW�޹W�|;�2]����$�Ѿj2�7������a�x���Dg\���rv����!^P�ɮ�|�7��ůX�� �(��dje��p���8& k���`�&�,���j����(�����9�"��E�#�f
^��5i�Oa�V�u>����_o`�X�vQV���?�b0B��`�l<�];�ߥ�b9�{����ʬ�x����{jj*��ɕ(T��\����N=���2vwv']�i�b�W�=��5���������G�HQ����lN��]�"�*M��x>�f\!�{���^V_���@�DMI�`�5D~-n.�M%���p|U__�<0������3
/�LMM��9��dN|�U�t��#��ؔ���bz��edd��ztA�G~��>�ğ�
ښ���8�-�K.̴���O�^��5�#>� �Q�OӒ'�'����Z�A��Ş�.4���������*T�[Z:�@=�x�8@̡MMMA���L}�K�\M�kz?[ �r��/����v��8�N�_RH^N�>��ؤ�����Xe�o �㊫/�*/��>c�A�*�mʺ� ۢ�{��WV�8���w�L<}��}M��P�w���S��p����?�D��l�VL��ծ��j OmLOv2�wt|�-H3�ͱ\�I_S�gD8��d!��
�S(sX@
D[��-��蝊'�Wm#���Lgg<"BH&O�GJs�r��<#�������|Qقd; IP���I���8�R���y+ů���*���#�����A�n�-It9�Λ��p�r��d��7����s�����.�#T�K�5���'J� ���M�W��!��� �3�Ձ(�&%���?T4���7 �[������V?JjM�k��fg�K�=��s��dC�/M�[��*?{�yY�:p�gV{b��x�7x�TY��K�B�W�W�)it��g�B.j�v��M5�'�r���A���@]��v]���9���Дk:R/u>���Ǐ�ϣOE 7 �A�={p���o%CNN�"Doe���0��Ҕ"ۘ�S= �^do�T��x��f�QIurm�{������͹uw���`���YۢF���a��ODۇ *��UIH,Н#��!�	R����zt�~Vx��#��I��7��-����Yc�OV+z�Ǔ9<6;;{�W6y�(0�>��KXدvp��-]�K���N���_�
R���������:Y�r����QD�Fc�:��CVE�#m(�������r��[�n/R�
�p��������D��j)����ڷ��C�����	؅� ^IS����c��rM�^Z�}'���ׯ7���J���/8]��G��9m*�R��T�E����"���l�=�_�h��Qq��K���p��K]�e���KC��M�}0�J�Gש++wss�hxx���~v@	����RI����:�Gl����'(��Bl�m�W�c4��1�5���vX	X��<ǅ�瀱��V�ՍP��w<�E� ��(�3���<�H�GY�f����gP���j/ahU+�.������ܓ���V�ȼ���5׷,���7��r��,��n�������vov�r�Ǧ�����JN�&1R�̑�AVc6| �feyN�]�\��5e�҆�G951>>y�/�eoXgV�ޓ�^`}1x&w��a��AK�y��鍄��"�>�*��Gú~�L{O����������8���s���'�^��a����r����@�27�7��pe�\W��\���A�i�-o#�N���K���"22ypQ�Յ����h��;�k%�T����;��q�>sp��uuk̭��-��`��r�:Jv�H����{G�FU�e�SS&e,�vs:�y�M=�"�ˀ�qj���w�����n5g�N��3Cy��GB2�p�+&c��p-��N��~˗���63�Ņ#]_�oe��X��EE�Ys�ށ�T0��/*����I8K4w4������+�{�Gv��6���9?t�B�`�oL��E`�5!!D�	�^�Ŷx`8�9��׹ݟN�`04mЊ�é2�SM�Tv�E�%:{�
���u!������cB2��vN��i�"����*J��K�o�k��0M�ɀ�%�5�K�'%�Y��2�/��8�5T�]Z�)�;����"B�aIW���NY����Q����Ft��o�i����B�͓���#�pi�PK�D�Q#����`��'K�x�'1Sy6�do1ۗ�X��.bbbK�W��΀a􀺂~�'NZr��ɨ�+p8�>�HW�2�� 	��j>���X�L����i|'�;2�3pR�g���@�)��I����6��X�p��o?p7��i��Q|Ǎ@X�/~�P1u�0SaT�iS{ �]\�M[XK�U�9|D�X�l�r%��%�P��6ϽɊ����!Q>Lబ��TP�x��Y�#G��m	B��Tϯ�ڹ�v;[[�����* ��.]�Ɣ���
���{��\}����Z^�9����	����q�%�˛����t%ܥ�\�1���4/7^leu�邥��K��)�xpyxx��� �!�����M��%���,��D��mX0��S"�$P|)����9"���O94ZddbF��@�/����eZz��w"d��['>�Tؑ"ӘJ�ݟq���ut���0 ��%��)��v��W_/�ns0;�G��'��
�`�%�@�)F�u�.9�C���\��J����5R7j���T����LT6���̗.G��Zz|�@����<LO�>�HaM=j��(��]��j~��z0�fO��r�}F����s&�w�aw�I��Ɉ/p��z��Z�ʣ0���~_tv� �?v�"t�1�.� �<uds�ч���^Q�����U�[DI�,]��� u�I�� ��d��1�qU��d��K��ɸ~.�����w��$��#z�'^�"U2���������8$�N&wt`��G��Tɏ���U.:�	�;�U�%-���/[r��Wp9]$/��"P��c�73���[�;e7bӊ����v�5itڈ݉c�r�<� 
������ozH��������GD��/4_��@�&5Ԩ��'Y�9֏"=;�1�\2!<t����k�c�����;�tA��AD�)���n�R��@�F�4u��&@�	�o����q�,�����}�.K��٣y�@��\d6Ms��*��b�З��?KיD�_t]*��������ML�O��A/�܃��8��$%m�}�Z��c�U�ǔB�I�qC�~���M�?==� �F�J���Wt�Xy��.�3
����E�$/��҂ک9��K���u��LF�#s��t<�^���z�9�����~�i�Έk���� +\{rA���$����@-��h�ª��4O�e�PR
Q��%
�a���S�[r�©�5��"΁�S�A��5���l���J��WP�Jl�w�"Z��q� �mqj��V+b�l�"b��;F�]�F�]Z�|^9��^��'|]W~r��������<,](��B��r���s���̃���-"����-�7������+��<�+��/W8�롿*SR��x��Cq�\�_���+6�j�&U�H����#����؃��?������./���cDxM��\@r��:�����,Z&%/~�
����pg�b�^����@�^���Ƹ�k�A�B�Y#[�i������IU@PE�'C� N�i�\1ZU�%ƹ�|w�`���]$�'}m�R<a�*������~_j6y OȨ2퍞+m�@<4��Ê�c-�,�� @�}�Lg��iV��m��Ŕ���]u��͵��Z�]}�+�DͨC�Xa;5�|�4t�,�fК\
����+cm\ %�	�!�J�Gg�������p���:zi�~�ONy����5�n��&i���;ݬ�����f�NW��?�]�z�`:�����!FH�DFF6�
l��M8�,�X!�'*����zq�E�BNV����t˄6��+G=��� g�ů��P�r+�mF��*��6�������WI�gS`�m=+9��>�sF���	�")0�y�|(���r �P9�29c�)QgC`"�J�˻��tXTl�r��d�¸n+�e�B�9��o��ּ������Dk��Rc7��q����g=�W�eX�*��_���?����+����2X�4BtK�a*����0��jy��|mY��Y����2�VQ�Z;X@����&Ͻ���HR�jZ\X�a�p5H ��CJ9�%^�h,f#P�y�VK�G�mm�C{��c"�1</`�1ZH7��V)v�6Uv��HrI�>_�}�KD<dm�k��S��:���������a����y~x%�оQM��Fh誢���C[[�JX�an��cn��a�V�� τ�sVJR�J���N�H��8�6�U[`�X���鏇���Ϸ�0�+�}�ZX�R��t�[@�8̶N�	��5�:���l��`�M|�sn�lh��D��
��0T8��xUP٬l�������t��O�dׯ�3��К�5��;���Xp�9��@k� �!�w'���+��"�Y+�Y���'9Hu�Y˷dv�q�w����u}��mr��_8J>L(���L�"�K���������t_=��KQ����jt�7��a��̬������+����ZF���Eh�V�aDQ�e�����7^}�Gxd�����g�0�A��I-QO�>�iS�3�4�Ghwvw� �.�D��VzX'?�G��n0Ie�b�'�2*�^^ ��nvQ�3ش��.,��c!h/u�w!u�^�K��~0V|jnnn��#n��S(ɴA����T��m���5��(�	KIM��`��_�9�^�;ݑr~E����]�F�����-����น�L)޳Q�e�os���u7  I(d<�+\���)orS5�y���W�§��!��T�P{�ߒ���th����h�������t[yl��!�rԊ0-[�fk�f�.[	���o�/�9�ţ��]�t��4rn������`\�C��ds��YV��-3e����ceآjv	ŵ�3�:0����x��i�#�'�],.;c�FVy�1G��+!�V_�.��ן�G���\R�d_
u_A��H^Jt?|�$e��������{%%��f����uuu���^2B�^Ԅ�xׯ_�mY����#ǃ?!��[J��DQ0v�Pғ45=��EQ��1��7��Ѕ>R��
�5�����X�,Z�������/ٛ���:&̣;$	Y4�[���W>��?�g��"Z�ėvg��i{{��'_�SÖ`�:��J .3��AZ¾z-�W�����v�[�c����@�{|�W�D(�-�f �S����f?U'�������Ը@��8=����� �Z)ua!�� 4{��2Y��]n�fp�q8lw��M�{�ȕ(������:�ހxD ��?�_��2�y��6��@l���6��l��qm�/ނz�HA���=���WW��M�&�E��7ۜ�-j�(r|�\�Ҁ������>����1 ��J]ⴍZ�]��k�%�XJ�%�,�vD��_����:l����"4��M���w�M�s�Y�u!hǁU/�Y���dǳ�B�ONX��}A�w�	�r����@�[��Y�&����,�Լ�n��VEl��%�3ü��φwcإ�S�E�M��Ϟ��{�;>::�/��lBB�"���*#;'�U�^�}~��$-��%��x����D
�"�]��X���Jy���=�v�5E蝘��	���o�~�	cRi|����Q�����Z�+����нg��D�M1�2�\��IB�-���{�H�M4��8p���;
x����7�0�8N:L�����6�u��tÓ/�w������'>�t��<ώ���x�A*C uP�vp��%�$�^;�t�.��:7v�������j�/��o�s����h#4́y3#�����M��Bn��A����0\I�.q��y ��ҞPИ�Vq�_��ԏ�i�����C*!oi���f�w�N��3)*)��3\��a5i�R����5�0��y����&~ߪ�u:�˭��\�cǞÁ�m����{?&���(�+w����P��QJ���w�㙑=�-��q�#��m`��+�W?��[9ڥ�%��-��{�k�Ў��km�+�fN��w	�A$	�P���i���g\�hXu!��D��p�DMk-jՄF���
[+��&�#?�,�Ց���7�2��vU=����]�h%�%�fѻ}9�;�rލ�/�oϻ��Bzc��]mq|v�]�_LG�>7�W��ٿh��'��J�n���ݔ�QA�;I|V�xF��(�F�чnn�|��&�;q�!yࣜ`�� BzRY鵠�|V�S�8�˦� �L�!�ӓa�#�efo���0ȸ��P[�i�"�Q�=���J�I·G�J���HW��p���r.l����������N���v!V��<��ܶO��2ao�ߟY��Z��T��I3��^9�dOf�r�n�����,p��,𱺱y���/�8��`':u��ղ畇���_�Q���Ż��fX:F=��2����B�.��5� 1�9�͖���҈	&&��!���q&ЃYC�LOߞ������t+j�U!h볺����O? ���4KrP�Dѥ댺z|8�R����I���55�+/?R��d;�^˚I�C��bz��:3��EP;�5���wЊ;�����mݔKk�'�S��ZB��
���0�Eָ�=U�� L ����߹�t��M�_�V�9b�H��_�0��JIs�W�u@�G���s���477��x8��{�EBB��5�I�Tf/�pm�,�w���pY�D���='��p5��F�o�;R$�J�GR�89�8�?u�5IZay> ����R3x�n����L�$��t�"ԳE�-sM��4�z@��'�A��_�k�BO�'տl齄�I��0ɉ*���X.$�쯽ظ�
ь�҈������ϧ��]>�;�ݻw�ǔ�4(3�h����$�,�QI�WW�b7,@a:4�l~;��Y{\�m�|�Vh��l	c;N=�-G�g���m������׍C�� �\�!���@�l]�gZ�MA.��mNNN?3��B8!�I�)�pf�K+�6�Lx�(G���ֵF�JG/��	R�H���~��4��-0�AA`���޷u��^�yr4��ӻ.�o���q!�LD[�`�=;G�B\�_ߤ2�)=��&�e�CW��qD��A�Rf�,����֍�d���i�$Mά�H�=~tbbb�c�ne0�EZ"%b�d(TM�v�wL�[{�zFi7ݲN�����Q� �ۇ������|F���� @��ʽ�O���V;Bk��ٹZ��ː��F�����j/����-1�d��|�%�gڣ�i�+^�3�J2o�^��I8��ne�8���L�J����e��B�91Z���F�������"~�k!xzjbw$3�!LڇV�qڍ�N+s��z�R`�c{�\v_�	.���q/
��X��d����f���#��^)���SB�����b�U��S� ���d(4������2xY &��~��8�c���Y�������1�E�K#(�p=+�U��������--j����j222M[,��ބVƫ��3E�2*j	�"̔Pe�
�p�ǩ8>A�@{�K	t��Q��QZ>+e�������Ql��#UϚ�� �}��s���>���uTB��˨(z�ɔ���v?y��A�����wĝ�|9@~�3I� ��+1v�>>S��I�x%��9p:�F��.�Ԩc:��P����҈1��W$4��K�qV��9���#/�ϼm>�(��6 �;�H���o��'_m�e����sF����F/=�E���w��/U���d�%�KV�w�p1@�T�I���d9�_����x�J�l_vߡ�]�b���D��*�S�����g�>�h'��l�}�u&e�7�����h�+7.���Es�{F�#>�E\!�DRV��3_/�D��%���n��ˠ5I���qɚ�R��t���~L�%p&3㾮~��HS4����r���V3ǝ[�<~��bԐ�~�8HV �;WiS���P��C�® T�#���!/6p|�Yf��UzkСV��6���l,Z��§ٺB~B>��Dˣ��%�5Cv�2#���Ҡ't�0���&�	�Ԁ�
���N�p�j����9?c��j�ٵ>$��)q3��"�S��Q�3���sK�K@�g�9�{##���9ù���k} ��-��� �Xq\.���p9��P{�����L�^ɌVњ���f,�]��<�]+�)T�z;��ڑvc�9�KݑO�B��%�m��\Ȟra�p�÷�	m"��{�����/���{O����M���.-��(�{��t_�{���K���#D�Bw>L�!V0 5�r����k:�����|�e@=�vww��������!h���iD���� <�Ah	uu�Z��Y�߯��{�|��`���j���&�clNh��?����L���Z��=v�y�'�B1w�IP�k�W:����ơ���`3��[0���+�~o���`���j�)� ��UϞ�oll���OB��Uk���o!�	uJ�>\?ߖ�w�GQeJ�	U�K���K��1ߐع������2F\�C��M�Al"��>�z����y��lv�ÿ��٤�0�r���p�G�������V�ӋTpn\��ii���'�4z斟��#��� [g�=�jp��49:�� S$��F��l<�~��nR2����n���1�N(�`1�Tkjax}3AGI��`����%�����y'bc��^?�(���Ȕ��/X�WBCb�9wy���s�%����9$��QV��f@&<���t%[�q=�b��q-�,�d&=���e�񝅘ZN����E���{���6
]_��Ʉw?}�tlfjJyqiI�%�h������
0V
�݄�]a�8�)^7���iу�zh�����$ÏI�Y>����ץ���9w�[w]��S�>�M*3xЛ˸|k��մ���ʉ��"{l��7_��_�x�#hM��p�w�plJ���X�yZ:���n���W9@��JE.��A�US[e�Gׄu�'�"�H�Nm�J�쪯���d�#r}}x�N��R�祖�o��Z�.��V���$0�J��_��Λ����X&��:?Ս-�����?y�a��y��!*H6�E8]O9;�3��Ֆ���]o�=�d"�`^�9�c;�7��@�6�L�ߘ��o\��A��a�c�Ԫu�\@�u��w4:����K>0Iwc����7i����n뀶����F��7� Y�ƪD��\�^� ��IN%�m�fE0=�y���t��P��szKz?z�R�g~gA&�z�����>	�9��i&�&��aco�Q���<�����T�L�k��	����� E��z�a"��2\�4U��p��$��p��:�O=�ᆪ��l/��R�̴�d�YRqE�Si`h��]�'�`Q%qAG5*pG��B�yΰfq��^><�.��C��K�K!Z�i}��м���	q��t��a�3&/da�h�{���n=Q<a��`]J�_U��k��
���CA�H����st8µ棖�73�.��<J�/��X���=]��D���le3���}�d�>��^*�ف��i�Bb�_�ٙ	C�l� ��eJ�W�(��mn����`pW�6}���ОX�Kzs�j��\�C
�\���J�X���ڝ|�h�Z\�U����]y9�(J'��p6�P��FK��s	�향���0��N���r��ba�2�N�>/�Wkd�9�� M-���a�N1_��&i{jζn8��m����E�op3f�v��禦��ʿr�HH�������|odV� V�fk384�[P�Bd��v�m~⦜��n8p����#�ZLP��K��U�&{�@ǣL�W1�f9]D�fE��w�X�an�������A�%"�I�|uk2߫S���Ȼ�λ����P�p����E��Y�q�r��JK��x&��vk��Cp��KP�J��*׾3���t���j-��8
pG������[-���V�p������8^�|aWKDx7��Ol�z�C��Fe���+�X##f�^��������8S��mɏ�@=~F#���I7,���#�
����b���n�>h=m���2��ֈ�l~]aD�Ƕ��3J��ȂT�K"a.�Lp"\VJ��"�ڙεQԣڅrz+z�,Ì��zF]v�SwF�n���r�{)���yj��a�(�e��0���;v�5�|�1A��<��(��s�Kj�#��?�����{���I���)\A-/��t���7��O"G)^�߬l1�Ѫ�PCI�F����������Lx%����D(D�gA�(�!�蒸y.ӧ]H,5����@�h�Eh��Nk�Y�^&�E[B��{���CU����3��b��0V�	'�/�3�	�c���G�4/űՎf�	 :k�����:������z+��e���0������R�� ����ԍC��A�Av��!�Fwd��o�w΁Pv��$�6�6R��K��Q��A
�z����yjR� ����9��[��!=�'��C������	wي�#;8�<��sF�Ŋ+-��p�S�)t�aN�;��{�fG1AQ�*�D�K`&���7{�����]L���/a��@�Z�* ��4��C��Q磛����Ӱ:1:Y'e�Z��V����ƫ=�C�n*�ƚ7�w�~��힗R\3Ҍ�th�b�y ��^����������k �3�yn��129Y�vDi��)�}ϣד�F����J��1z 5������bӔF���2����)�I�ѶD�?�wm	I�f�m����A��㳋!@j�f/GN�{��dlP�;��<�l(�K}Jd��O�R*�[;3�VU�p-�-u�	fGʲ/ޅen�!�3x�o��|#�e�`ל��3�������:��g�N���/��>b^9xۤ��ܵ��>�W=:{�i8��r�G��E�� [[��ǰR�[����/��e�-���Ke"�k�z�;C.{d�v3��%c�=��J����RJ�B��#Tg�D�����rе,uY t8���,��!nʡ���4�Ƚ[�D�4H&RDVX�L~Y�=��av߾�E�@�mJ�"���\�G��9O:P/�
�,o�.�W�=*� �
�ä�����ǍaX����߬\a�K�~���� ��]��`����kU}V�x������	�.}u�T1=*6,�](�l9:�����@��xR� ���&��>;�~N*טe���8���@�1�H������8w,��MJm��#v:Y{\�K��� E^��w*��lW��C���k!vj�3�E-�1"���F��N�ׇW�f1���y��t���`G�g*�V6�����;U?���*} �������H"Hf��:�V��b�B��NΣ��Gz&[��8?v��;��EH����&��n�6��1��ԃ��c����еҤ�M��x
(��N��)t}7*��a��)���s"q�Y�,�+Q��</59J�"���a�/Y��ʥ�-�bF��3�eU��u�e��W�3���v�����F���y��/3&F�1�.;� u&��i��X����] ����!?�N�s�j|��	�w!�p�m��M�3�c�t��A��{Hބ�<,8�&���/7�5)�mZA����Te0z��3��xw�٧.��v�cj3Vb�Fb��n:��)=jnc��+�Pj�������]S��4Ҩ'�.Ru�;	5{�k�֦��Z�#�0�����#x��Q�O�(�?<��w��߼4��K(1.S���������k�%�jH��a-]D5���S��O �w�-����w�\�@�̯�9�W>��Y"`	�8����0�(����ɦ���a�	玦��C5kph�e�K|)����9@�XH�=`��[�c��=����Ws�,��K���z�G��C�H�`�La�+=�Khw�����>;����Ʒ�P���+	:TCN���i�ͱ�쳎5	۵��gfL
���7 �L�k�3%�Ŵ�9��Uf�1�5R[q$���P�m_�m�|�1�N��"��n��w<��/�}xxy�d1Y����O��`x�g̒8��6K\�'k��۩��0fJ<��w�o+-;����] ��}��o�����ށU��q�˝ʮ�:	�����.�����;��MQ\�������7q��b^o��}Gamn��@������r�X$Y���K��^������f��;�My6^G�Rh����0 ]:
�ĮL���Y�Q��v.�T�L��.�$C�>
qy��O��U�v
}�8^O�gH��ed/��	�h*�7R�L�G�;�X[�B�-��wR�l0M��	y���nu�Xo	9��-�lၚ��JS��х�GFvF2-�t ^0h�^��GC�U�L�m��xr �wl_��{�&="BOe� 2Ę)9�6�R|���H�ͺe���ڍ��'���BY����q�#�py�R�0�P�n�f��B��<v}Aǜ�!�,���u0t��H���f��ȱ��a�MY�l �E^����jx�l��:�RE�48��>��n��q~{�R����o����O������3�IPQ�����X�8�J��=t��0��� �:��u�2���J��a2��2�/"�3�,'��Кx�_��qj�e��ޥ�#��Q�y�B}��{U�}�]@h��C�6��ǎ����z.����O(�۔.f���'8B.�i��{I/q��o�{�~���c�C���x�f�Ceqv�b��՝<)����Q8�	�q�]xHf�"��ސW��V ��.y;�p�#;z��K)>�e���/�{C��Oo'�3��H�s8	��bڵ��&�X��u�4�o4A���>�pW�-{X��m���<�)�`
^3��'�G�S*sHy,C��HG�_�(�:�sa������pܺ�z�VylS�*gB�d�a}������2Ό ��&/�H�٧P���׉4K�g�͔>!�"N8 �s�p,�����;nhܙ�LƔY[ ,�Lח�uI���kG#f���531=�fC!棓���و1}����$Dx� ��������vh����넌x�7��ۖ��	����_<{�os�~���������E�q�D�E��DR���B�k0����e��E�5�� Ǝ�N}܋�_$���B>,|�@"����h�l�'�� pV%�{���W�"���K��9�I���H@�*�/��%��IG����H`���?���k�d~����D����}�*M���PK   {c�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   {c�X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   {c�X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   '_�XF&�!    /   images/aa671e02-30c2-45f8-acb2-14f46084a715.png��PNG

   IHDR   d   (   x_C   	pHYs  b�  b�<2�   tEXtSoftware www.inkscape.org��<  �IDATx��[	t\Wy�޼�wI3�,Y�%y����=!N�Ҕ�@Yþ�@��ۡ,'
(phiI�B
	�,l	Y��N�cǋ$[�dY�H�h���w�{��Hr�=�=\{4o޼w߽��}��c��kU44M���'�j�ڝUT+���������^�Tas���ɇ�]C,_����R	6���Kv��h��׼��x�"���Bk0,Ǖ�@5�Mtd�WD���(s���|<�`S��6�����*ʕUzWͩ�d�T��o�8�r	�NM"/£�f������9�e܍��舆�v�".y�L
sM����<�6�D6��n��8�U
��{�.�|>T��5ݎR����
���f�[�Ē��bĢ�r:�TH!d���9"�7�V�A��¶�!�z�P8���ũX�փ��f�r�g�bGE!m!7ڃ��
�v;�J �q`C��3S(����� B��~|'q�=w�vJ��"����c|���lN����}���e!�����H�.HaC�'&sx��V�=�������J�jr2B�EY���,�g4�x���h��J��躆���r�)umc��Y�F�����c�M�R�M��Ahʦ�KY�h6mU�۴e+g?<���D��ʰkeL�C.�EI�hw�#^tb� O&VxQI���Ɇ>p�:_q8�y�KI���ྜྷ���Cb��?S!l6����$���߹i�z���4e!N�o������y?���֗���!�.���!�/���|� ��R\T�`�!�����f���xd�l	99��+��D�\	��&�>�]��s��8u�^;S���R$E_Z����v���+eԷb��d��_ن�~�=H����Gvߌ{㽈�X��ē���N%Q�W��lw�en
�z{\^�p}��ʕ�jZ����)���~�llCFa��g��C������/��JMȗe�Rgoc�X�T8U*����)�R��a(�m��C�2��L)�R�2ƿ��w?>���K*�\�=*�?%�s�����x�E/�/�g����i5�t.��+�p�x��8q˔(v4G�b��|��c� )��(�W仂r�2΄x�C�d�!�!���2h��6���e���7ee��?����H�((.͍!37���Eo���놌�]]����y���4k$F5(Q�o��U�q�m*<�d �^����#�;hL6[<5�ΫdK���C9w�ǲh]c�A1��X�E������??���o�F���Wu�I�A��xW�+�JE<�lF<ځ��)���s�Kn��A&�2��JX1��]�ӋiL	4#��5�ʂ8|Ϊ�lˍ�U�A�t�eMi
��K��_K?�~��ى��s!L�9W��C(�k��ta9�Rr�ƾ|}J�����,�N"��ڜ���P�,�q���t+O��nE�9I��U��-���r��t�^r-���÷8_�uV���W`�D���s��%��Ĩ�~\%Z������Ԅ�E/��4�A�
�%���G�Ђ~��\��Fx���]yň���B�|���x�jZm�e�Ǎ�[�oL�얹�m��F�G%4���h&v�Ӂx���ہ�&��bY�m���J���:���߂͏�)��d�?���t�J��������pߊI�(K�W�?�7��b�$P)v�J��o�v��w�@*FΑ�U�eX��^���,e��\���<���R��xs����xow�Oy����<��RV�?йC�I��m�����M��,~|�����pud�EbI8l�`���o��aA+�P�\�����=3�}�x����������9����ۿC�+b����A3���+D�g�~�ʋ�06���̪<�6�
8L��	J+!�++%POk���F��o���x���!1�ο��q�bT��j��y�s��A|��sQ��h�y�4�G�'���u�m�M(e4�F=K,~��12q.���{a+	�v�����6^�c�V5xBO����־��'6�H)��( ޷uc�i���\X4�q��e�Td�����v�I���b��1��s(���$RL$/�ExeAe^�3t5��*���ma8�N<u���;�حrqE�[X��%7|B�]4�ʁ��r˚϶+��Π
�%�E��P�����X�[�R0��	��D�g��V	�6<3����N"�+��U��#8>�Ɓ�Zh�Xv�Ex��$�li�=O��Z���2*!{���r��&���)K���w�a��y�K7�c�� �F�W��0���v?�=���o�,�L%�Q=�m��^E�	�.,�6��񂳺�wd�d�qQ�[�mEH��t�����ozu��m���]#;� b�C��6����c52����\�o�H��3�>���56�q[�$QqY�L���܁��_�A�zZT2ط��5�P�F�ǰ����7Q`II��h��5)�8ω�)C�2���?���Η����q9�RF�幃�B4�9��W�丢cx6�8��ɸ
VTa�\�q���6��7�T�O��]�зi���"��E=౽��~
[XW!��^�έ�I�vU�2�nU����B]���^7
(p�.�j$y���9���s۱�ţ�+{Ԅ8�M~|�W�+��NJ`� ��^
����w���o����q����G�����R�G����Ŝ�� �~�"��d�6��cGwX�\�KP��LJ1�M�5/y��Sh�GW%Mq������WF��|���q�p�K^S�-,|tKSeB�k���
��Cm�h�ގT|���a�E��	_0�2!ʨt}ZsG��]؉C�I�f�y��Ds"��!�� 
��ꪳ[�2�ˤF廌$v)�OK�WY^�w�E�?�ǧ,��ŭ�pL,��݇��w��qَ(^�{�T:J&O����vpz!'B/���"�`QP�S�:��#���e�$�y_�$�(&2Fq��f|9I�;\�ގ��A���B.����������?}�ե񝑵�'�*�Й����p���R?:$I��Z����c,t��C箉�:~`��&uwCR%<|h~ER����O��M�U�g��=�W̻�k�F�hk2�07����}e�O���xB}��ߌ�B�ED:?{�&cYl����*��[��Y6y��p�CbxL�?��#7x� ��Ղ#�x��r�>�O�㫮��}$1��}��n������e]�q��!~���|x}^e�|�/J⃟��}aD:�V߬��1{\���n��z�ۈ�?S
��H��bh�G��ݶ����K���g�"g�3�]T��f�#�o4s�T�ݶiR)csi�Qh���2�nd�Ud� �q�Exۋ���s��z�>��ݡ*�,�|8�\%+Z����+�CYց*���R!?̌���mp�=�~�a��>|� ���{��ij�<���,�b������;3��L��ϖ����ZH3�56��n�>����S����`[V�zVd�s+��tw�s���gdC�~ 6�^���ۛQ�d���W���h4҃c����O�������O~�������{qe�.��z_5P(�r�%J�B��~�"��%�A6����:�o�+�Y���^�%��(�sJ(�L��*-�jb����=	/6�o� �BP��D^6����h��^ANEU4�e[Be-A'�Kn�U�\��p�'�b�a	���D����B���C��:?�Ų��<�~�@6��T��\H#�/�N����Ai8,�fr�T\Nˣ�2�hȋ���q���������5/{6���\����/������"=�}�Nv�����l��Yxͩ�a��l�e�R��Y���pɂ���x(t�Y��0�	�K�`�u�uc�MbZIA�>�Md�Is�cr>��TA�v��x�s��k�TQр�����Y�k7J"�cB:9w��5�%QsB�O�j�R>'���h��ʠ���,~��^��|a���BL)��M=H�O�u��XE��y�~�P^w�V|��'�-(���a�FSLL��zH��KHrOIL�Ġۍ|&_�Fd���o$E�|�_�f�'̜�E����;�Ea	�
�E�G!�s8�rÚ����u\b�D���]�G29%ON�6�l�<kJJ/���s
b~AVY%�&>;]D}	�^�U�2�+���+77����8KE�y���<�kU$S���/o���k�؜�뾵��=!����{�w��c�9�$��k���~7ԏP8P�ɱ�8��'в�ê�b�l@`kD-���l
�R֜(tza0?#��C$CG+��˪.L�
b#�g�8�!��@O��*�00�{�xì=��G�� �v.�S�wl*��HJf5/,�̏fːˏ�bŌ
��S�I���gjƿ��x�^Qc�������sNq�������,�[I�����lƩ���?�5��)�8���2��w���g��"Ǒ4W�&a kǆ��HƬ�c
�|��-Te�ԯBX�UR�lϞL.�A`X2���)AY|W�̌%\�	,y��(�M��B{n3���?:�E4�R�9:�X1��|ȹx��u[)<.�%�2���<� a��'Yi���r�ӉC(]��ׂ�%��ᮔRa��r�VHF�j���B�!-h�c�ZT���ju͐al�����^#Q�϶�?[�3�w&xP���1��/%�qۃv����vy���� ���`Fo��Q�m�+_�
��v8]nu��^��ϋf�rW�d�W�z_prK�)�q���B[y2�H�VT�+�ڻ��2��@�q�UW&k����#bqDE<��Ev��F���a�nai�01�D�|d���5�A�c�b.�
�V�d٤IP�B�R�=�KƐ��R}L�/?3��+�V(�6�UW��&�#b[^=�ࢋ�F��K��O_����YMVW/����3C'�>t+���-g��b�(.�~׷�X�\�;�������k!�{CxD�u�
�bU]Qc��|E��`��&���B1��`��$o�`����nlI!:
���j.�F�)�&
�5�R*js�R�<����R����Z����\��_\ʋB�I)Cao@���'�%��{6���Or�xJ)-֩���Ǧ�/.J8�v�[1t�kTaQ��Q�*��"�#��U��V�?�`l~S�=��J���0�s����p"�����y�[�(kK����b��[�BYDh�>BY�3�ד>��(��������bC>Yq|\s�Y̫�&�����ěox8�ǰ�݃��r&/�oy��[\ʩ5��d1ּ�,:����W����n\r���Ó󯻲�8�)i��g7������h��ԉ��X8�O�S�'�h��j��\⎓ʺd�VOp;4U����!�,��zU�J�'t����k�S��x���č�B�@�!�:a/C	�jSU���1d)���2#�3I��x&2|���:���m���2��o�AQ�m�i�OZ�{t�`��pv��(/�T���Z�

S����;�?�O{����v���~Qt��/�~��mh���8���%ƛ�G���k�N�c*�%'�����e�fNY.�Na�1���^PB#��gc	Զ��N럊�B��?����pʗ�!�|H*IYT��u��T.���7҅$����;V�2��&�`��|聉E�q|QW}c?�b)�K.r�;:��e���]�gdZr���� ~r��V�B(kl�d(;�(.
݇O}�RUl,ˀw�e�U�e������-]kj�ڥB��)~R������q������eȝ�wg�(����C!��l��א2%�����U�d^�K�(��w�Q���uv�*�dב��;������jwesĂ���ϕB��|<8!1?]W�#۔$4y/��IjZB�����.�sx������Zs�Us�dhm��3����
���n�R̈́���Z�ʺ�RD��,"i%��v!k����z�d|�SD]1��5R�;���Kv��KBse%t0>��WU�3)��>���N���.��DoK--���3�QY����F�`����0������C�n	�0�!����G\����91������7BW�sk֮�p�0E���\6�VEU%Aq�_�~�dB��-��Y'���eX�ξ�R
� ��"ب�6��"d$���ߞ7��\��<tr^�ۻ��@u��8.C'V���=/� ����0�O���t�woEh���{xa]�)���v�@�ԕ+fu�*�:	[S�X�Dfn�rzBpx�
S \�"�dlg��Be���*�ֻ�j#���k�կ��<'�dQy%w�̘�iA`�˪29�1�lmcj�6���H�˵}�:����!-���'T�h-$��=��rV�VC�^FUľ�%������A�L�a�C��*�!f�^q�x���it��b�̀�a�3�^�O̧���[U�Ya�tOMbt1��cs��߮���܂&��i�ы�@�|&w0
��s�"�LkeY��#1���.$:�Y��+�U�ʫ�@^E�
��p���>W[Sۛ<ʺYBo�d���I�^G�c!7֫���ښa]v�o�`���饄�E��
�^�{�{ў�DE#�p ���$�e1��W`C+�˿���	���f�:��>&Qe3���8��|�ׇ�%Z�h��z�A���J|�_��������&c��\7z�4n�um�{���Q˪*�[Q�0V2�P���K[�`�T9���~��0��
�}������2����[��E��|�"G����*��9L��0��ᩔ*8��{,q��28T}h7��J�*��֌�ebsr��4�_������^�Z�Ru
���ƻq@&5]x7���۰{gQ7�Ne��� �;��pd�'�K���8��Fx뷔@��&n����E'2g�#6G+�:<��B%������B[��ϛ;HXza���F��G��N/<8�Tװ���%��R%�bņ�g/���5c��¡��1�IG/�Z)�
ɠ�J(��zQ�*pWBH���t�v�7��L��Et���|�����\��w���T���4S����Q�Le��2a	�/J�{��um���΀�	a�d��	7m����Se������A��B3yKm�X����9�(ֲ(x&x�>��h�Z}L��|����.^��!��2p[��\�
�O�,fʹ���s1�yX>��*��%�c���4\�3�+Y��f��n)�5!��D����3W�dW�.�o�H�7�~tZmAP��TC<������2�\-T��Jyrt^��w�S��~+��-���c�;�{�de��b�;�vr]�Xߑ?{���X_ɻN��ŵtc=���Y,#��1��1����߸&2K ��&���A2pE-w)_l���C*�T��L�w�B8���S��ڌUAqkw&RYL>���ƅ��?$Z���X�y��fZ���bx<�.1��4҅��s����E~��63    IEND�B`�PK   '_�X����?  [G  /   images/c05be033-d934-4815-858b-3a150ff9d8b3.png�w\�]�/����B�&   54�(��- ����R)�A��N�	(J��JH� !�@Ȇ��v������߽w���>O��9s�̙�Μ��D_���f-�G���'��;K�΄ɡ]�?״�c`�;~��BڹG��������������:1��yy�9<{�$��뒵����p�A��}���ՙ�l���e�nc�S�Q��N��~Z�M�,N����>,��ہ7�n��Iӛd��b�>�[��ዎ�տ{/��3���J���s��]8:=w����]�02Q�+�Ȅ*�(�(㼣��2s��A6@xF\���o�~	��i������j'/��8���pR�N9���x|�q��~������������|�_���og�Q�_X�e����ր��<s�A����S:[Q����b��O��
X��T�6�+���E,0�!���{�j$�J���,'��p gUM�Q��5���fTR�1Lf[C"S��1	��ӌ�;?+��G�����
)�e����y�S2ۡBp�/��di-ep�y�<8=���ʩ?�k�|�����
Jӗ�V6O8O��㧀�!�&��!Ì�!�xly2�"�g��ʿ�B��~��U�����-)�4�p�A��8 ���f�kԅ����,�����}5[$氡���x �eRl��D2��Œc���s�u�2�Ox��M��Dj�4��;�ۈ�F�$���]cl6Uǐ��ŵ�L��_�푇���Nѡ�P�w|s�	��bC��Os��s2���y|�����X���z�|�)��~��۔�+� �
�q�q��dv�ݽ��Ț���v��d����x���k��^�(�O��z���	|{��l&]1��۶������vL��U?ل	3Ԅ�q�_�O�p����}GLZ��
�9&w�FM�h��������T��M�vX�Q�����#ӸF��v�?������2����O�Jo�+b�//�Y�{�h~��vgjkA�)�g��Δ4���x~jF�������k�OˍO��v�oH�mh���ϧ�l�XF0nw�������n6�=���d�4���	�;�r��Zc;��tMT'g�V��� ���:y�h��cd��ëɃ8v��G��Jv3���]�0�Z��:Py>��7�`�#90�CB����E�F`t��/�+!듪�Zr`���F\�򹪙��y �2�� ��SX�!�N�i��F�V%pZ���l�����&z�T�:�$�TlJ���|#{F���Ư0����k޽g�oX~���&?�7��_�H���_�cY7
���������֖���$���
�A�bB��XN�L��ڂ"1��^Y���z,�}lT�ڝLS���{q����-�K��@�p� :�*��X饸�����X�k: ��j���!�z+��qT�q�Y�߯W�6�U�oi:����v＼������ �&�?�v�k2g�OT�oj�+ *�#B�>Dr(/��]���N��ʶ%�/s*��C�D6�n7_d[aD|��8+�RD\�:�|�(�O�b00��N�K2�W/��5U���LݮKF4��X��o<꯺OW7� �����ڶ�I�W�T�5�<��S�����T}7��Gu(�^�������(ڨ�[���ap�|�9�h�$�-�0D_�J.����\��T�Rs?�!@q8GG�܌�4Ý��(lـNPx�v;kwXm-���k"�N7<�y�(
h��;�[����n��#���A���8�{E��/�� �m ��\`C�<>�E�|7���n��@�NU�n6rEJ��d���A�HY�m�4��fhjI�H�_�5���	G�;Ym˿����X?��6�3������bY������������'.�V�6O�ҥ=�}�^�JH�xᢩ��`���;�/r�~:} �SȀ�ϓ����Dz`Kv��䉈5� ��1������h�qs�Gk��L1c��HZ��g���y^v�Қ���hW�I�"��|0}�i�&D7�f���mcF��
Ǎ�Ѧ����_R�����_�O��􁦁�І�n*o��V��1�6F�-Z���|-(��[D���L�h�۞4��_�e�&�-�
,/}�_�юTk�S�V���ϟ?yHR�碣\>��ʛ�R �9�q���u��+���&� ]����5窟=|+;��O��-�b��^\����/'P3�����ܫ%��gBl�Q[����f'P�[R����ۃ8�d�����tl0O�1<�X"��Ү�䒭�&�\�A�7����T!��k�tu}��bs��X$�(\t1�n���E�s?)(/NV�9+�B}-~�'�ѽOr�]&U[���#�7Ԓml>^�-�1R�l\�_�G� &���m�ņ�������������R���E_i�0z��t�=
�j��.��m���@C��>?\թMĭw	(.Uy�M�W#������&ؾ櫧l���e����T���bU�l��q3�}�������3=8���L�z�����7�����/}5-h�����R�i7��dQ�`��~�C������������)
෭x���!���V����T�ƶև]�/�c���cԏ%�W��!d�,������`P��֬�#Z�Y*�]>33�B_��o,���5��v6ڸ���p��顅hҧ��a�h��ĩx�Rn�ê�|:�*�'�]
|ҿ���#e�Β����9�����V��s���k)c�����`$��M���Ud��ԇ����e�93�m^I�S(i��AS�V��������Lp3�����.���K�6B���ݹ���M�D���
�'��LՀk��7Am2�3�Y���f~�����{\?��@;���ίL��q��b�/��
/y�Z}h_} l'�	�u���Jxrg��<,yp-Çu�
��9J�!�����8��R��l)(++�]�Tt9@�1+ta+#������ M��__37J*,5�pm!W�� ��M�O���٩qppBm��2�������5|��a�2Q���.��/Ʈ��8��U-��̓��Uy�l7o5�j#y{�
�׽�]8C[��B}6踟mN%�"�����f�8A�S�#��iQ��0V�aק9�jD`5�ȯW� ۜ��,�F\�r����t$0�1c�dKf��g�B�߾$��o������T�<�G{ş��`���!��|;\�������-Z�?�m����`H~�`}�7�nz�`C�C�޾�U����7.1aww�H�~� �]\I]"V`j��5�f
U7I(��q�ߗ���|ىI`=��X��7]FcD�pP�6`f�4��β��ڊ|�j�g��]�хe&�Ω���6(�w$�I�W`��g�T��]�
c�3ۭo��߻��E��GTt�x�hyi��#c��f%�;o9�2E��GO�^�^��Q����h�e�YSUvu��d�������'W�)m*T���
f�\�<�?1�]ï��곺m��R���ߑ���"����T\�vk�Ό�L}N҄��Ϛ�5W�\*���g��Ъ�P��ofsp�K���b��~ŋ��B�Al���x�H&���?̹����zv#�as+�����Xl��Ƞ�L�fl���	&f����;����_m����+j�U\��z.r���냊t{��Q�ūJZ��l�2ޙ{�*K0��N��c�o2�F������î�����}�ΌR��ښ�>���O~��i�F-u��d��s;_�i�*7����0m�W�(3-�vP!R}�:�'��];�D����|�I�*Iq�K��W�E�!?��6��v�FZ��m,��E�2�[���8H��&�!��}O���S+��W��G�S\����U��VHi����_��X� p7�(6ല.�2�m������4�������1�K^���ʒVf~y�I�"u ��D=\���.��+%� Ga;�^��r*��Ҿ�'���s���u�oc�J�J�ugO���Ě�J�����np+�oDs���lw��+��PK�+�C�8���hx�� g��d�)�{pD��_Ƙ�0'�)�z��R�J�%%{�|e+8���6ǿ�m��d��=���/����L���> [���N�!�C/������/ӫ�=��36�h�r���w��ǽ���s�s��|Br7>�u�B�!.)�	�ڟ�P�P;����Q�n6�{�(x��a< �-��W���}�3\�۫���H1��|�̚eN
�	Z�m��'v6g��K`�3��l���/q���ޟ�����/4'�䱥��E����d���N�a��hs�L��U�H��p�ĤQ�vx������Z��^�ÂF���~�]�RLa�_4�!�埣'��?��sO�)�4,�����ܪR�h	+��o���z5��{DG��0�[�vG_��7j[�E�����0�V�������L�Ay�����ư��c7K�&�OHg-�}�}i����-�v�[Y��Q�e5bt��e���6n�3����`�ӫ2�����ޡ���5�T���Ǆv���%?Un5i��҂��3��x��x��˞(-��Պb5���q��Al�O~�ٟ�g����^~��!�3*��n���z�ȯm�P��O��}�l�x�뾯�[�5m��V��Uq6P.9:�/�w�3R*S��ll� 9���芆�ш����Ko���C
���`E���g������i��è�X�!����TN�op{2W-�ln%_Y�<�.6�81/�����r�W[OI'.�?
?���`ri]@*��Tf޷��vf�cq:��2�N%��r�O/`�s`~��C����(�BvS�1�k�3҉����V4����n�96}�y��#h��<���`m�MO������1�|n���G�4Լ���/5��-�V�%g�p�(���q�����}�3��^����*Ї���vcqu��7ω�s���^՟}�o$K���o��˖��y�����4tFP���A\5a�o�>���K�h`�z%���l�=f ��|�f�l��P��v��Q�P�:
�t�xL���&&SI��C��f�ܛ�g�]ޘ������r8�`%/���,��?�@�ݪ)�U�@<"ou�����|�Հ9c�G��L�ʒ��{�UA3�U%��9����E�d������;q���[�Q����")B)�P����[����<3������}Ve���H��+���m�=�Cr��Q����t�Z1�����5	S��2�u�R����]5���<��l.<(���ؙ�r􃇯j��'�s�^���f���5����΃������5r����y�6�yo	.��O�o����' vEﮍ A�I�|f�+���L�I�ir�P����/�cu��5��<�զ_�8+%;��k�8m�j.��ԇs�%gDzF�v��}�����~U�.U���w`�b�MJ���9��#"�j|VsC?j�'Oph��#d��OZ�k��~���"F�z�I��nO�Cay}� eS������w���܋�af�h����mr�^�k^�͡ߣ'�ȵ���E��%+r�~ߘ�GM��t�E�CX�̫�s73	�G-.N2Đ���f]L�Gb�J��7A�K{�3��ށ6V��_�=Z=�"6��Y����y��ޓ@"����de\V:����	F]�V?��VVm�==�����χɅ�x� r��mqō�p���g?��7��f���x�W@E��4�QRIW��<d��s��������sf.'\�m<�I`X���d�7h�u�ݲ�Џ��7mϵ���d�tD�y��B@�� ��UB���̪��x��鮴M̧�+5-?�WӰZ���z�/^+ ��'�=Ό��~��wk0C�Rׇ��]%����a��/̎6}v�}��
�r5 �Lp���;t\���1�V�����)V�����:�B�fS��G�� ���1��\1�gZ�^�X�i��.D���۰���d{s��7��3���O�S<�4�|I��(�NiwV�N�5\�ڹA�{έ���x+����p�?�0�,P��ă��Wv�'2��rY���&�#��!ئ����7�-����R��Y7�m�!U����Bx��H[��M"�E�X�6��v4�vd��+J__O�`]�ycf[9���<XM��GӰ0�#���B�_A-�EE5��������K����#�P��qo��/X�]��f3��Y0;�r#DG��B�8в��� ��n=�e`�7�}�����8��L#[r�Y�y"V?��'��Ȓ�� Ő)�L��&��#�p�*�\�<	-s��z�lN#����]���
���Dч��Dpn�О��N晧`Օ��>|ժ�0^�T�
�Re����	;��I��Tl&�9���KQ�!��.�@I3&ؖ�Z�6�MÍgexq3h�MI�y��Y���u�?oc^k����X��8���˝�m����Y!�fW����>Iv�< Oé%K�_����*��5k��ޗ|�TQ@9MAa'f(������O�_FuY��i؋�'l��f9/�M-��E|�) %0����7�%�^&{��#Ԧ�"��*\?~��0{D��Ʊ�+T��J�]n^/P����������a	��;2��A?@sqg�w}���E\΃�tb�q3��ң��� �W�_�K�	�)v���g�<�O��kX��ޞ{��H���lK)!�A1`΃��%�~b��a�r(�#{d�A��vNw=>	iJY��6[r��0y�Z��36��� �0�r�K`�����n��ER���j�^�p�<��0�6�N|�y��tE/E���,-}����i���N�e߅�^��7��}�2Jp�mM�[��\B-�< ؘᩫ�%ѹ0��uދ�W~���f�n��NDǭWy���2wGl� �U,��ݍ��S�"���P��E���cp�����23(�p�j�꟦�ʹrɛL��rƭ���-ȦR!���[H��t����~�ăS] �`�@��[�-�k�B��.��X��&�x񸽃`[��{e|m@��p��vaO1�Q��h�w)0��{ҕ�N@g��pY_�{�qY���S�����hn\E�h}�>��;��˖U�/^���M���9N��&�O��:�/�N�L׵�4V����|��\㬂��:h'����C��hxcvT�ߋ���
��2�D�&��,�w&Q�Fv���-�V�a�����;�0�?��X�ͫ�^$'Q!��K�ׯ����9lM�LzdI(3G�dv�V�P��̝X�K�so�/��!l�N�5����"h�9����&2����JNS��Y!K�����r���?Ձ<�>��H�����piA��k�9��i����>����e^6z"]�,�|�o��n (��ڏ�?�=��Ӳ���|eU���[�ᴙ��@9����܅��'G�`w�����Q-�\D�{�m���ْk�5]���#X�ԍKϠ� O�y�vl�R��3�>k�u~�>�%w)��k��~���:��UϖW��\><��1����2,�fWR��Ө�����#�s�� /��*ʯ�x���hsa�F�l�(Hĥ����H���?��s��DKߪ�a�W�[툣�����%Z�,|R	�����ƚ}�(������a��i�JL'�<�G�Db�k�~W�Ί���e��۾�زQ�0WȻe~)D5�+˰�Gx�E]�,4���b�˟`r�����g�b)J����|ޛ8�%s�ecY��φ�\��Y%r�>�ݯXyZ����7�n,�6�ᕐ���������ReE-	%f��ok�f}�V'��M�j�M!{c�J���Wj��rKh�����߬�`�����"j�/?��9���韺k�k
�<��/��ݡ��[~��M_#��K?Xy��X��D|����.����>@����aB��9�E�Yx"kK�t�P�#oJq ��'�<�72O[ ��};�����Ȁ��o׬��ՙ���F��?��u�P-��ǟ�0����U���r�����)0$����9ք���-���5�4Y=�F��p���7
`�j��4Vz�e|��m�.�U|�ʺ��i�M�)�H�{O�"�]F�9�˺�,��:�%T,�;���:�`�p++��#ĬC�%�P�?�L��q���7�, >��?KɵwJF�G�������Fy�G*7����=�����粌�l���G����T��sF��3�����W���a �W���|!�)�֍�g7��#8�ۖ���'����Yo�<=}�>���$��T_n�'�憠;������~~���+e19-�?X�a�'�/�W����������	��-Fv�ۋ\ъU@��g�5'���U��2L*y��Q��fk=�R�n�VKadH��$��<�X�K�^(^�{TN�l�O�Yo�i(�l�=[ƭJ1��/����A�<k��!���wg�Z\� W�[�=2����ӓ��3������%.z�xx��w/J�K����9��Hמ��/+��	T��,�Ҿ�-I�{��e��ͨ�L�znB�W�(��ʺ����<@X)�^���ʉ�]̹���x��.�L��X�LtQ�R��������3�u�MI5iX/��uZ��V��6��u�U��s�$4�e�$��`p�����9��\��J��DQ����0)?(�	�dw؎a�<pU=��?�b|�V
�37�djߟs`|��#鞷#iwa;���ndG�P���z���x���zuV�BT�bu�T'�g�@L��$j'�"/����X`�L���)>�5{��Rv�#j;�ztΡ*��b(F���K��b%=.��T��Z�L���S�b����w:[/�w����d�6e:�׉����R�B�9��<IA����~�AgA�:¯8�/<�͉T�!]�hz���^�8L#ll�m�§+~�(,�:`�.>��@�\R��U�V�O|�-�y�d�=)�B�.q�ȹ���[�A���H��Rҽ;@�q|� ����n��x���� n�Xk�_�-��u킝��N�A�rw�\ �/��敏_u��e7#}`)���-+����@������$#�ԕ��,<�����'Tߕw���u��k:���}�����\�}8�0Ll�@�"�a���a�1�����嫧���&����u���mI4���G�Sˬ�鏓~y��"r���=|ex��������?>|n�ݤ
�OwM�lb��'��x1�.�;Uѐy{�	m�bC��S�-3\H����TιD�}/:�+�/���T�WvEڞ&�����Ν�e$2|�����M���t���ʺXC�r���.�\���<SVaɇ��YO�,˙D�*��}��q%'l�ږhR�F�80�a���q*s�t�G�yٍ�$��N%�Pw����A��7�����z`H�QJ|�ك�oSWiC�Iw0�-O��L<<�z/����3�}��hAJ��
\_ܮ33�1"��!Z�a�T���;����0d�ZY�����3�.s��G�(���ط��j�m���:s�P�MG����d&p:�u��WedM���f簎����U��裍�����b}f�}s�m�ٷx݈������5ՙ&�yL8M#���8�������Sq�8�P��w^,ߕk�XM�I�tW��
K�as�����y��QG
��Nt��pȤ7ޖy��Q�l%Q�l�Ÿ�=E]X��sfx�k#l�݈,�p�;m�@��KN�0�2�Pl�U��h	��������\��x�6s�H��M|���r��0S ��B�����Yٸ�d�ct�<����gK�z�����1��H�aK=�����"�����L�@^��v�ZZc�(��MM�j=�0�mÝx�>���� r����K��^V�u^� H ��J�r��
���W�����7�x����P��5�[����7f���#W�vqia�ɡ-R�Q6����#���Ѝ۝�M�w�b{�%���v�f�k�dq��[x����׈J�e�����>##&�����"k�ŵ�*OU�}�P�lcX�!'��Pw�B��G=FK��xCh�2�m��N	��T��b��?�-g�R#�-$�l<`Pz�d��<�W��Fܸ�'�#+e�6�-i$d�[�<	�w�sA���2����|, �ѷ����
1L�s���-o���0��	�^8�TƆ���[KQ�-n/_}"FHGĄ�I�-}x�՟���	N�f)6I�	::"�=�j��;���t�:h�\J��3��\PJ�mSU���O{�z
d�T��C�+'-NZ������:��r�Dy�H5���x��M�{Љ�D���Ͻ�5g�>~,�\���$��%�IO�P�sw��b曲���Q���c��PE��p�@pel�#�&D�1:��*���a�wQ��Lm�sH������Z�!����X{�M�JngE�����`*,�8����yw�c�VrC���;���bE9X��#i̴�x�?,C��	�$X;L�~0��RL��m����=�c�J�	^}�����@�� ]f���@s���o����Q�Ys��V.���R���������]x�ω�;�B�R,\�H��|��}ʱ�q�>D/܂�u�1GXJ�4�"��d�*�~=�Q`C;a�z��7���~0..[�v�ƻ_�P�PRR�sK�j�M����	�M���^[�J�) A��������I%Ay�M#~��Y�pIY�p:j�̗�<׻����#�B�W�^�������ٜ�~�zG^E��ad1"��O6�cv�L��ަ��"Y!-�WT������+4��%|쾘�}�wu���]��D&���V����1fDǷS�{6�����b��J.�����1������nQ��y ز�J���`�bЍ��?�;�>1r'3�i�	�4����Q�Mw?G��7)�)��@B�+EEyT�%K��D]�,)j��%Z,D��*��\k>]�� G�6��1�TČ#	��f<1���5+)�V]]�on�(o.�QQb]��J_gק_3��|�8�Ɇq���$�?Q��4�Q)�}��(���=��^j���]0�IY>���}D�K��b��%4���M���|4�V�~t�̾yh?�����:�|e�q�z��R��e���(imi�������Z<y��	�%���n�Rk�z��C���r�
:̵~��yz�c�gӺ|�ϙ��
�2㟐!�����X����%�ѝ���:���6{7��o�ם�oU$�yƚ�e��Q�r�N���9%�&�@y�kI߃F����R�_A�Ɲ^Y.���;X�P��s�_c�]k���EU��!'�u��م �I2�T�&i��TWJ���X�Q}��o=<�:�i��8�+Ԕ�����"Q��Б�z�׻��﫿���Q{��t���:Z�ʤ\��r�����^x=�.'���D�ޅI�+��8@���ٺ�^m�b�ӝް�%�V��]�^�s����Z���g��ßN@/��� ������W��؅�c4�!p�.���fk���UH=�=����y��jM�ȹ�::{���r+��r�����IIz�M�Ka��|��FP��D�g���ЎMn&LՃ�����o�\R��zY���c��GvI|D�.d_KV:��]����g�	�ʱ�
;��e\�s�8�<sΖ����#)%8H��U�~Okb��9�'С���1E�Iĩ����^0j�_F���m�=��z�yrMe]��s��1����SW�a�
@x�U{'�������28OIbd.�;��G:�PчJ��,'p�5'�����.�6p����̠y&�� ���lO]��C9��Ek����{�H2�:�]>�pj*�"�[�r!�#��0�=�9����9ntͷ�}[7��m�8�3�k��c�=�_r�Au�{�~'S&��WLP,렷�d?�L��9���$�Z�eA������5'��pt��s��u�Cd)�C{��DH4}ھ�gHʕї�H�{SE��Ʊ�����WL�*��ϼOC�X�����pW�pl���b'�厌Kt����:��O�v-�������?�Pj����a�6�dKM4b�@��ӿ����b�|@���V�NqӵD�>�12V#`�;Os�ߦ�zI ��5T}��=;{e������E /�`�jV.>S����(n
���_�<%t�=�)]_�)������w�p�ԇ�{+�~5��M�vh?��l��/�ŋbh�5R�?!>X>'��[�v^�����u%z���;�,�Lu0�g�@�;~�ϩ凄��&�w�te��r9��z{�*I*{����!bν]@�(招�����a8��[�Sp�Q�d�=��o��`>������e>y;N�z�R3q>|�����~)�Y!q��n����E�,(���&;j� ��~��E���m2����5�|�&M���+r �W���]�J�)��=^I��8l]���˺����ѡP���1�3uD�$�KL�O���$wd
q*����1���ꆈ��������(�p�RR?�!�F��G������('��O�$ߒZu��{�6�iY�����6R
��ft�I_�� �>�mi��Ԙ�����Eu�A����ȋ!.�[��N�W#�#�et�?I:p��T��Ӿ 8�Co�i��6�}-�O�?gf�SRBOo?��5���6��7ԍ�I� ��}���;WM��D%L��LU�8��U�
��<Ȍ�T�^v��(��#=o�*�-���S�"^IY �1�Ig�
�Y^>�}�в>`{�O� I�&�t^%+�G�~×.�P}a\�r�ے�\wmc ��yN���z)�n=�&2/3�,�����Ɏ��ر�G)}�;�����V:!E��}����u��e��hF�t�9�g��*����>O᧥��k�]{Y���b� Kh��A��v���Ğ
~�:�ړ��:*�%�0����gRG�+u$��W��VT�[-�
:lD�=�>_r��Y����Y<IR}�Ӵ�Ra�e:��<Q��� ��ZN�}=�}҅�	��0K���Ug親8x6h��3���?�W�kV���	���Q���W�S�,��Va#�L�Ie�@�'�3�D�&;�;{7�޸G���~�Ho�_���q2q����K�v��-�*|y����E�f�1d�������^y��Uf���,���/q_����d?���+�����
0�F:�[�O��oso�����>)���nڹ��@y~��<i%�+��4�U��(��q��\�U_ ;_6ߋ�\��E�6?��Xg���͠A7�$i�ޞ �ZA!v3���||օǚ�WH8pJAn	}�z=�tX�{�q��TY^Y).��<�'I�6��z�E[H��M^;I�7W����yKZ*_��@8�+�����7W�,kj��]�B^�,�o�s�4�K��3%ջ�:��.���X�Sv��6}��?����#�-�g���K���/Y_��}��PVZ*LS����>��z�r�۷��Z��o�wہMj̍����TV|FXN��E��ӥ?8�j{Ŧ]���C7�K]����N_N�P~I8�K����K�R���/���O��e.Հ�SWK찥C��b�ɽ����tqth�.�i�o6`[��~8�ߓ��q0�'$�������̗���
/��i���$�-8�\� w�_�����奡	��Ѯx�?�.}g+l�@�=�=p����ZX��V���Yb$=2ݩ���^�dT,�ɼ�ۜQ�]�<^�{�.�q���o˵T�v9�����)3���i�Jz���3ww�����l�%����iz=w2G���ʟs�j���x}!�{��h�]�	�%%���FFF��=�<V�C��?'+DR�9�؞~\��*�����
"��/(�H1���&{�&��0=���W5=�59c�ʮ���]z�m�L�˳&�}^�����<Yd]������E[��Lt�L��z"`�r�<���>�zeU��Q (!�f	ڢk�.K-x)�T~��8�fo�^�e�?6�M��R+1�c+Tcb;�Α�g����E��������⧘���� �*r�dr`@�:+�[�ǖ�#s;��p��<L�	9�me���_�q���E~�������#���U�<����,~k���R��;����S&�Τ��w�K��4��޽̓���*������@@��w���q��E,�����O�5��co�5$S/n�Фy�/'8^�-T�/�N�]����r�fl����G��+|4w�s���u�a��y�+$���M�pw�LF�����GY�Y��c���C�'�������ր��%]|||&Mhd�鶡�@.tn!Z�%[�o���h?��/w���hO�G�xڲƾ��V��i^�s<R}kC�Ջ��F[k�^�I"qO�Ύ�pb%lt�")����V���N*��C0��uJGo�[�C�y�-U�ևYbC���R�<�q倅'�E��,�Vb�Ј�΅��uI��f�!��8�w��;ſ1�lY	�=C���2�RÓYh\����6*���>�LG���14麇Pc��Vk'�y7�JI��v�C�H�+���/��S�xg��2��dq��,O�H��d��(V���7شN��oF�L����r�R)�:)���1��܈2f�A�=�(e|�#���$�Z������M��w�A7��9��#�K� !�o�A�=�f�|�+6��\�jI/=���aC�#�R�ԅf�>C-�x2X`���]�)�x&f�c��A�f��P�aF����%�G���d2���Aƕ� .�9���0��0�[��O�W8��8�Qk�u�H�ċK�b'��~�x�V	d��	�8��O�%����CŻ�����Zu��?&��X9:Ԫ�&�E	���V}뾉+,k	�by��u�c(��6���N�mI�-���ILYX�!h���e�������c�y��u����_���!�0ic�B4�I�Ξ	~�a�X=[.�8��nO!�U�I�r��[�b	���Ѷ���_Ðȧ�<7����k��V�s���l���W�Į6%vYu�FB6%=� P��cs�qc�ю�ߣ��ƌ�c� 	;c�+�[�X�E��;ӑձ~bw@���~�u4�r���[�z�ue:������z�<)fM���-���d���H���CCk������' �z���B�r��jC!]]G�O�h�*λ���5/�7*S������#���|�u����Z�{=��o#@b�V���>�
"���mg�;�$�]�ײ�����:9�B։�n"DۺS,��Y��^�����G.���"�jW��r��V�L��@0���HD���(�(R�̃�k��ŽF2��7��F�!���^+r�эM.�c���Ճ8chU
�&���7!����+%:�Đж�@\��e���B�ʽ��l'��D��;F؄"���M�o��"�B`7>Z8E+]9(�b�ËE��f#E����5\2�x�V1����P�H/�,E�^r@B��̆���q�=��h=�J��[���Uce�5+X�Ɏ�%��
��Tyܖ��9�'5�����k/�8��L���e��W��9P=�픅��o�h=G�݅`����v^�l��Ţ�.&�̈́��&��f+4A"w����daU4�Fv'�"����d�_K���[rPȴ����~�g��7�Q{��2���k2��5�(@s�ܠ(4З�O�a?N^���k.��#"��g!cr�����?��x�{���JӶ���M��Z�����+H=���hs����|Uނ ��d]�(X���Ϧ�;�O<V"n��}^`_USEdFh���Wj�Y4���5H�K/8N2�{��)�߯��$�4�4�0th�4��n6p`�K)��-�R����Hԓ�q�ՙI�����c�G��^�/PK   {c�X���لO  �� /   images/cd9a76b9-8a14-4d7e-9261-140514b5ac3d.png�XS��7��*�QP��E�&EQz�Ì�( HWiCE:!0E���;�H�� !��)����y������޹������Y{����k�$�o�)m�rp�6嫗488��98�m���|��g���ʷ7�?�M���檎=��5�o�/p���p���➝	�}leno|��D���4�(w���0��n;GN�t�&w�M��?���\�^d�[ox�-�M�3Q��7�o�v��j���
'�S|�BjyI��00�m�5@/�$]{^�!��J�WW��o������3��~5�X����n�x�N�Xc�n�+���!�Y�[�ĩY|��/����(��NsHG/�ȤyxԆq�%�b2�R2vZ7�kR�u=�כV�Y�
;�����a=r��/�|ߑו�����Mkڃ?�o��.�Խ�;|���,����*���5B�ؖ7r&�E��nZz�������e��g��6}�bq���j�QRR2�k~[3�lM��Y��-,�_6m�h�q��U:?��v,
�H���1���&\��n�}�s�ti��]�vij^�	ٵ뵉ά�b1��D1繄���+z[�g����a�g�J�7_V�T��R3>��Y���qΉ�q�&0�������}wwy�H�]�j�ς�կ`�b�=73�c�yR�a�g����3�����~�τ�,J�f�hPt_�5�{ .������A������^�2���,+ϲ��k�i������N�p�ixy%�����XSl(���^"7/�������677���:.���;��������K.$RUS��ۚ9c���|�ϩD��K��n%v�OU��47��@'�3�A%���X	F�!�D�������(cOOE���}4��E�PQ�٦/z�#m`;C��r�*���Z�XP��*˄���OEbF�@ �.L��-�EJ��o�e.�c��JN��6��b�����~��+������l�&:��F��ͷ)���Z�?+���o�,�2-�/��Q����:Z�e7h>����Мf�����P�X|aH5�y~�J�����C�Ζ�jA���b��^ד�.����v�Ym�ȯlm�މ�M�(}UD�U�I��m��ͽS���>�����
�)bi�?"l���\&&&.�m�^#Ą�~7����S�P������2-�agC#��f���2q��I�ɡ��55oj���t�b<�p��f|��Ǟz:!�bO>�dp�z.]���YS���V_��\�c��X���#sY"����sCλ
Mu�Ė�|q��	�̗��(jX����d���m׹(��^4rj�#;'a�+�D��ͽ���2N���S��S�C4�JV���+ɹ͋{Щ}U����,ݾ��DA��"R	���k���2��Xn���N���;�:Ŷ�wBjy	�XE&`��[SP�rL��i��U�`7���7`�Mhpٕ�sY���P��l^y� �D�p|���Pfv���{VVm��L&�X6�h��}TKK����f�Sb���͡�H6Ťyqy�ciD��y�����n��׬�p�&�%�?I�Mf.4�z�ϒ���N�����(l�%Kd���������{�oii����TMg���y9��(�raH>��F��8�0�V5I׏�1��ك��}���C1�s:r��(.���Oc䅔U���g�X�]NUC�_�OG�_M�L�q�Ilz�דF0���w�g2�'��7^N?֞)����������!#��(A��]�y̺�,���o;te�O�|����(>&��v��q�W·q�F{w�{��B�?�4�=Ļ�e���fg���㭜��ǘË��[���®3f�޷+%�Ŕ3�Дv��w���գ��]tO*�:�aSa#YK`.v���U|�F�d��@9���y����kJ�H-���î�������\�if^���%W�ܗ��!����˃����w�C,U�.�7��/�4QI����dd�l��)��~���6�Ɋ,��4��$�2U�m����>2�Y��lf��t�iCtE�,bt���+�^��a�P��`�(���;���a
����0yF������j��>��f�����5����}�#���y��鱆ŀ�<k���<wi�:�v%99��LT�3a*��`�:�Ƥ-�q�x����?e%���-��`�Uh#���S���EEE��[YR�[��Տξ�˳�;���#���|�%V��X������D&�XU�4I{��:�8[�ܤqE�Kt��\���.��Š����/�,��a*��|�1��
-M��BG��������	op��CS�
������(���2��5bw����ğqB�G�P�f	3��%KӵaL�]v9[
prrb�j�����9!��?���$&ɣ��Z�����s�Y ���`{d���/�/�z^DEE�WgV�]��2�	+��}��������������Gnb�˞��)`�e�߉ZY'�5����m�W��Y�NnS�%{�����mF-���{�5��i@1���Ӹ�,���+ڃ�GVVV"�ԋ��K����,�)B#��=L9�S��A�6��v[�\s�<�:!�<�1���j��d�z+����/*T�[zr2H���}�Hi�2u���(���x��`�vS�.)4X"�2��
����v1��^gW�KK;���,%ŬY���u�M�7�џ=�\��]@�0�����g�H�؛��i�9x�~ȳfw��y�}���0���f���1t�B4+�r��|MBTZN.u�܏M�����`�07+0-{�6���YN�Dd�!)����	�e��A��A��p7ڞm{2�@����wt<�
����zbO�Ts�$�A���H���k���,�F�1*���{�x�[�u�o��6et}���O�rm?k"�����yK\�y)w��ň:ט�b���=L��l?g|`�50+�":������l�l��i)���p�؞�`����bf���VKz��w��~���KN�p�E��i�r��U�_��P{���,�D����9��gj�S@���vUv��}�8P1��<�h��]��80	�g��w�/1�e�M�
9���.{�"�����,�F<Ɣ�����'㒓ۻ�Tn��'�����dgE�66w^�x|brR�jąː�R`�6d�'�C��I�xiŔ����8���i4�b�AP�ϩ2�]س��O�dؼuH8���+,��,��L6�e���3�ˠ8�P� �vo��~�]S`.W�x�b#��]]IA���򗰨(>
3dK_���T���X��ʦG8k&�u+�6]��dP:�k��E:?9yx��V����ٷVTz�Viب�[#eU�UlR���F;�������ƥ�3�l�}V�Ŏ]QG$RSs-�L+�����D^+j���.��s�B�sخ�cW��3���tu?�{w�v����|�"cbl���M ��'�\.�ɺ�|e-+�}Yּ� I�|��nK@��6B�UֲU����ԏ9x��v�����Du�p�ɧ�1�{?� FI��y��/�ck촢��{AWX��_O�ð�\�=)hVΩ1�aǆ�8��j+��Jr[β���+%���^�	^^�m)�-��Ω2m*����GGo�]�2��wE�P���R��VMO]��`�j�{�#��!�׏��,��?A�6�1�O�#+���	ۚ��1���?���7����47ֱ=�ڲ�G����=�K�kV�\e���"��[�#0bl��e�}m�#.��Ҩ�*��A��4|w~�;�V�����Y�草͏��l��Odk���T�G�TV�@�Y�9F$���@�0,��N�H3o֮���I�6!&��(ё�}l����x`z ^�{y~$�bS�'�����ǿS�V)�/4�ܡ�?8�q������_�����ej��5e�q���Yu�!���L�Ql�\69�ᵍ�'�{�������f��:��0�-�NA��\O���x��0/t�.�f)w���j"QVb���@@a�f7�<g#��s%���s6$�b���셜}���Ma�H��"��'8��EVy��%Q�]�9h�r��FMx򨯟�_8��^��,����|��S��M�مOkY3�%�k�
u��/4���y`*٫�^6��6No���3Od��������:���'Ϩy�������h3���54T/��D�+���ND��qt^N��J����d����y]9Q�e�����Z'��--O�_�"[E�	��^��Z���
�raV�q*�� ��6�S�hY���l6�W`w���Ȫb���ۛ�x7���ҕ�N�����z���i>��^����L�������,Je|ݾ+���\3v�zy����5�	�]��9%�҂����.��d�nd��xKR�V�Yy��:�T�s,;�!��ʦ!KD��Z�J-1h�pE�=�,�i�W���,Q�d*�����LP��!��^�C��#�Y�Ȼ++d�,��:I�BL������6�W�<�h�t�4p��N���$P�����B�������%��qI�r4�{�b�M+b�W�q�S�V��g�Vb�r	JԠX��*����a�M�Y���f�%��	�ZY�����`w,
Ov=�Z�<N�*cc�es�☕Q��S�����ρ����g��\�z���\N�"�]��Q� ��m�pִ[�E��b����2ƾ�3��N���T��/�*Dy&ᾣ+��!F]��@>R�u0�޾:��Rk�is]箳頕F��H����d��N�弮��G:�B&'q�Q�iii�=û�o���W��"��Q�6Kd��1]������a�?���daGDD(�2�]���Gͼ.U����'���V:Ű�6K�����uL_�Z�^mq�H�}q�$�a���Y��[,�����'�}]J�ۧ��#��o3j���\��N�/�� O@����x��+�`��ҋD�S������^5���'@�_'���Sw� 8HA����4g�������{M!�$��(�V�hmְ=��xlc���W�����:�b@8c�Q�C�N����8w�Ձ�a��N�Q�U^�[zI)q(��2FG��(�q&�)f+���z��C�de�/wP���~PM�>׾bnn��Dg���EU�*�������'е}z��Wؓ�g��U�tt�a�L��7u�q��˛�Z;K{H��}@z�^�b2U�Q�R���Tɣ��Մt��?���sp���F��d0ga�vB�yy�6�u�ۘK�"�K�j��2#�fN�f[��^$�U���c�J�A�仒ǯw��F�m��>����Þ��?ZsW��Z�������������a�C��Q�NEG(�I�خ�z��E2�qb~^���V.��
 	V?��P�%Hד(-I�l';sV���уȑ%K���M�\&�j!��6�ȃC��jUU�����a�Q���EN��D"�n PR�$��O������^�	�h����~?��e�hr[n��U�)��|�#�hJ��=���-k��y��4�Xw�=ü�
�f\�$�f;4'��&��_$Y�>�8�>�@׼9i;=\�]�#�CmԤ���<#�X��1l�T(�D�.�C8����#��^�XQ�~�B��c�v�X!�o�����D�� ����F,�c���TJ�@�jVW�o�cQ�	`���N�1�!:�d���G��%E$4�?UVVfzH��_�MT��f� �f2�z�X+h�d��D�>���L+���W�͚�
`d�?�Ō9���N�l�ߧi�63/q~8H���зAG؃2��0V"���	���d�;�����
�Y�������K�hV�|mV��K"���_d̩h�Z8��o\ܣg0��QE���E����0|m��Ս��42���E�����+��ݰ�2L-f��6��ӽR�Fw�*�Y:H�������3W�r��84y�����ئ?%)*�;x��-�^�^�'ƈ�c��*8��ހ4:,"Ԋa�^;ۓk�w%4��bF��5ms��M�n�y��U�	]g�I�	y��f��5����4�|8��u�))1�.3:��Z��b���	3^.��
���H_�u��Ը�6��H��l�
�|��򣳺��K`3����"H�S#�w8���2��P��Z�!P T4���4=t�sw�1��0]�� A�M#�P��3ǈ������ޠ@M���"�b<ӳ���#;����;Rf�|���GR�?��],A�Br3�m����D��$�Kg��K%��7t'k�f���܊?�SKP%$��`��e�"E��Jqϱ,j�@'_Ŗ���n�F���Ά{�w ���9���O�����F��)�4��z��'����N�w�U�u���ʌlN��3_J`��{��D+�u���_.��Z�K��H39��ܒ(���B���d�B!�~�ub-B���"#˰$��@���,>����Nv7��p�NNs?}"Zv\�Tm�;�T�8���+jA��_�"�eF7ݦ.�@�A���GPn>˝����D455��D6�m͵tԧ�}�K�,�!�HGB[�
��������o
\�f�f�n���,��j'�J��5�fT0���������&IGy���'�0�6�j$���lOk'����uY�H���Ƣ��r-5[/5��~O=��I�y��xy�qWng.z�e#^ʼ72Ƽ�f�=�b
��d��ׯ��<������������}�}���o��6�ovQ���b�0Ϻ�?�i�W@�����`e%���۾}��ĄE�ъ
��q�i�L�"��r��$�Nq3�a�ё�8 m��BLCaz�^�U+I1��Mw�e��cO�}����ǂ��=��$3Ɉ4�TJ�����(Yį�L�O+�H�B�+��]����)��bZ�w>���I��q��ϊ��}������LX˃3I`�ł�����-y�_+�L��tC��js�+k7�Zy�P����*Ǚ��2rr��St���������sp��7Q�+�f�އu�I�;�&&&�Aj�l(B�P��#����_r��W<��k�v����[��� ��6D˧$�Ǵ55��@3�rPV�&u''&Z���W�3ؒ��򖓛{�8�ted�[���I3l[XXHVZR�	���֔saׁOn�!ӘaT��9��ٲ�x���RS�ua��<����4��vvUUU'}{�r����� !H]!	��B+�&����e�X�r

\�: 3>lu�2ڕ����N���KF�ZH"S��^������r�T�_nc��m��#�����eeS:,��,,긕�:�NǚSr-S���Wb�*p,Mg��֘�����V�F�V��d��1^?�ztf�c��V=�s�#8��������@x <����@x <�} �*��y��u:/��p���N�gz`#�F�N4�Jݶ�,�_I/�F0��`#�F0���g���OF�[���U�*�z�#�F0��`#�F0��`#��G���W��+��F&:3���'���q����_�#�F0��`#�F0��`#�m�}��*Ϧ_oR�y��uod*�o�������V�Oi
��i���>��j�/�^�A��?���c��W����U��a��@X ,��a�m�v��K+������a��@X���yy��r��������8�0^�g����X;R]��C%�"�+�����'��G�J^+��Dj����'�=ڹ����N=��WS9~���ШqᲺ��W??�ͱ�܍��A��j��瘇S�NY�]<ߌ�W��?Ç�.rK�rt��\76N(���ҊE�C���RE=n�3��Y�С�!�Gq1ٕ6������P�TDm�UR�B<��|b�������bm��W�Kt��Ε�{��?vX$<Ohnn.3�8<���9��T�hLD>��a벯^���!�C���ώ��I;��ȗ�k�ߙ�$�XI�r~�%�$,�kr���2X�O4r����	n���%�,�k�!�g��C�������a��@X ,����lfٗV�`#3�$62���ӯ0w��+b�[=0�,Fb&�\!�8���s�_�1ەv�=�N}��b2!�I�9GN�#K�O@߿w�Ǻ�◽J�=�V˺����M�L�w���+PC�V�a�T��s�CN=&�w�����:9�I�)�0d$��4����:wb���Vzv3��g��Le�����Z�PDQj�p6�0T��Ɓ����`�b�
L1G���	��+(�]�L��']���T�sP{�0��� �ǻW}�����,�w�U�ȩ���{���w�?<�}��ѭ��	
/��P�l���uO�������?�����9�:d�v�IߠN����@X ,���@rҋ��g���a��@X ,�'�-���B����$i9J~]��(&�'�>z�W�ڬ�h�uV[�`�2O�jh�zj���W��yG�ʝ�)��_U<���e�"1R��"�8��F�,{�,M/���sj'{P��Kxj�u������v.s۽��.��C2M�B��E��T�ù�����l�F3�2�V	l'E��-Z`�	9޴�YiO���À�%��=�(�F�(����Z�b�C)b;�v~S6�Rҧ�ɜ@6�>_���?������z�~���,��/{�@X ,��a�����",�n�\�9�-w����oD�|��ݛ�З�y�����.�c��x��V�a���� ��`7O���.�[z+�M�׾O�H�5ڻ��~�Z���r��+��r	���r�������o�wp8[bh��z�i�wv��*/bES/�9����'н_��fc/:�㻛J�x����;N,�����6t����)iF����@�QKl�8���2@;�D�r��Yh�+G����x��~��)�ӫ����X ,���7:�ĻC���
��a������_����-�`#�F0��`#�F0��`�c�70.9�ԍ�l������[�F0��`��&Jx�i	}௢�`#�F0�����O�|\��N�EW�nb\���F0��`#�F0��`#�F0���N�ڌk�W�Y��J�nf�~�F0�[#��کU���F0��`#�F0��`#�+х�R2�e��2��`#�F0��`#�F�A��fH�Y���^0����_A��&�wR�F0��`#�F0��`#�����KɌ~��`&�`#�F0��������m���E��`#�F0�ۢ��ʸ~��N
#�F0��`#�F0��`#�}Q�y�Zƥ�RZbf����7�wv���`�?��-]V=��F0��`#�F0��`#}G�qj��۩��zt�MP>i��Yڃ��#*q��յ/�x�4#�~�/g�f	�%Y�W���3��s�`b�`���G�2?����L�������������!7c6Z/װ��2V�x����&�:�~)�~]|��u�z+?�:c���L�0����j��a�s�gjۺ���;�?�`@�@�IO�W�E���7�	������6��عť�Ԓ��8�Ϣ54�M�cS��:)������r�{��!)��p��y�76ځ�$�h�Թ-^M��j���*�W���7���������kybJ<۾�+Xz�I,��c�v�-�����5������y�8rG뭠�]V����Fn	K���7
{k����� +���f	���o7���ܑԹ�k*|O~��:95�o�B|Zåޞ�G��hqe;�&7��q8E�����޲�ߪ�����j���c�p���r���U����"�

��8	z�e5y���b��7�R���������o�ȅ���`���dZ����y�7'������by-��@F*�<��P��
���\+�[ȵ��C�л� �ˊBu�7��;�b�Na�Ah]kX+��o�"۶S����?8�\�L5�Dr~cP����H��P��N`��	`���i�s�7��S�}��ޛ�am�� �]�>1S%�m�$�ڋ�ϭ�����zt��z�|�����[P�Ruν�uJK�_�����7��c��^�f����W���h��y␹XǑ�΋^2�N�mP��1N*��/��B�s�	�]Y	s[�Q]��+��r��2F[�ۀ��8��	!Ae�bs�JUߟ\�aؿ}�Da���dg��b���1�^����m}�!,���u��lǚq<�մX�7��'F��1�\*:L��|�cS���k�]p]�&��x(��|Xk�g~L��s�̠5��7@��0렘Wl�q������_�ud������'��ˡ�a��^�V�V�V��)����fA���T�0^����P�sUd�"���Vk�}m2���呺+Z�y�/sآ���
��O�x^�*�,e�E���^�q P��{"�JЅ·��mF}r�}Vb(����k�LE-IQs�'.\lK��FZ��A4=�M%�G8�'��2�f����wQ)��Bzo�9��6���u��ha�$C�����Rt��Ķ�p
i(yWf��m)�e�	�٣�'z��*���ߝϖ�-�����:`��~q�YX����:�NW"8�{��c�=�[�9�kZ�FQo]K����R����ʴE��¹��~�0dw̦Ϟ�>�~gcB��:��	H�2!�o���N�5�첢��b�p�G��g���C��C��ЕA�g��u͘[c߯��^=��xBM�i�f�e�_9=G�m���������˃t�vR��<Ց�%�C�[�H���.z�2y��"{��		�6�k 77f�/�h�8�����N�:��<UB����ܞ<�m��	�)��i�t�c<�<�,fmÝ������.�hz�\�<�[���}<����י��2��R�ב��;3����R�%��s����o6]8#�Ӏ�+��q�%#u�4m<�	rQ8��-�m���+*-z3~4\�V]�5k�6�݇m���y
&���`x]]�[��	,:�p�p�V�`�����!)�"�p�t_���_N�7�oT3�ϐVK vV�t!N=�yh,=���zب#"j'�`sYa>�F�F��ҷu��3������ƥx�'�n�h	*��'�^�o˰붙�m/R0\XT�
�C0WC���U�h����@�[��K��D:����(ؐj��_"vddF�-��Yh*��i���5`ĵ���s���F�wc���5�p�n{�J�z��F�t���Z]������r���'��+�F���k�@9��j��h�)�q�G�/����k?D�7�@��X�*����-a6�Ԁ�y`p��o�����uWHDo��D3���k_B�t�9Ɠ���&�m]�=h������3��8����_o��)�D��f.�qyr�e���3�#[L�B�(���ي�i}.�=���)�8��C��-Ϳ
�=��%;������t��o�ܲ�}���^�f��y��DҖ�����@y���缓�����X�0���ȶ��H����H��w�:�\��.*���/~3;#R?��X(I?����=�qX�����R�|Y�ZJ�� ��]饌%���i}1�=�e����rsþ.Ϲgf3Cg�Q<5�u6gf�BRi���ͳu��#$S����Я��^�������8s�)n�K�rJfD�`�;�t7����oA.��.on��|�GJ���x���շ���VT��8���1ZYf����ڬ㉷hCET/�����o|H�$ta��#�7t6��hC�$��;��ť�4
���y����b������z���û\�w�� ��a�O,�LY@�83Z��v��=��v�?4fg��帞@<A���]4\���\�4�Rt��+�A�4��%e��|u���/{ژ<���),\
L�R���=/��O�]��SH�� A�>�^��c�]��*�G�+���<U.Ut���é����[�`��'Ԗ�Vψ�٫��[��쒥�p���Q�H󱡁K��w�4�K���h�t�h	���Z��9W��d����'���9!/o8���{�'Ч��m���#p��u4��������Z�P�fh A��~dxH��;U�Q?�*�*wB��Q�������<�~yB5��uS�ξ��Q�RA����\��PQ��P;�F�>��cP/�S��w���qo�n��܍��/��'v܆D��
�������V2&���ލ�����}ת�U���^��ܪ�ڗkKw���:B�$�*���wb�E�c�=��e�z�*g+���������Z�Z���sV��%*:zy�gO��'����\��˪����N��[r�k;-��n�� ��҆��n�V�n^u ��*�	�>H����gl>}�^���w��|
=�5�P���t��������K啯!l�>A�Bܥ�ң�	5),	�A�pwV�1*�NW(84}3�����>U�+Kt��/P8��_Ҝ�z�hχ����z�� 7R��g*K�q���G��|]�Cx�|�辨��bc+�O�������@;�C�m��� 6Zx+k�yd6@���ّv9o�w{7��s)G0@t�2�Nd̤��������~��;
E�N�@��ᾦ�׎���V.�jҪ���oVpٗ�3Y�>E�#���a�F/4ħ�]����Ju�F��y#&:����v�8aKMAi����
����M�-]T�+aȲ���Z�{!a^z�V� Qa��y�b�P����T�)�	THlo�����}��e7*!72�f]�Ŷ�ȗ;WG{S�����sA�?�R�7����C:x�ߣ�vэ �煥�޳K�o�zF�j�Bn>2���/w�h\K�ߨ�<�D���a����I�Cz�I��v
$����>����K_��m蚾d�賠��0124�R�6pc%E���VM̎�(���8ꄦ@���[���'�@�C���h�x<%��׸����C�h�����?����_��X�1�Ȩ�_�]�� S���!U	��Rt��ρC��R����ȅ&��<�B+@l�������%A�������1�.{Q��@K�^���x�KK�6NO�dD�����B��W�:��
�Y��x���z5� �I�f��~�k���ۺ��竹b� w�2�mf�����JX��p���S��]>`�"�õ
C�8���y|M����kJtf���Ly����F����'<ύ�C(x¨yB�����_�@wT�B�G��X�R�m��Z0�Tĉ�q�zh	s�VH/��"K$��+w3�qi�}��Q��GwM�N��9~�T:B�Ae��$ϊ����x��Zuϐ4.��kB��Ӈ*��W�4�(�L�n��F7���S|1<�'�ۺQ����WW�@�-n�CO�(��-\�2�͈�昫�_� �cTfppv&�V@f�Խ�R�]Rab5ŽBј��6u�C���Aq}�e�j7�lȲ �Z�������K�ڐ�@�V�C�f�=?��D�3������� ���O��������2Z������W����+�E0�5K�
l>��W�aK-�V��l0@��	583+�ae���O�z��fM�OB�I��� !i_�cuR�r?Ŝ�;>I΁��T�	m3�i���R����9��'����^�PX
�Fk�Ʈ-xw�B	�6���15#A��=+T@��,��ǽ+���YO���h�s�U�b<�d �V�N��P4�X��[��5�DOnT�{0y����	���x����
�%�9���yB��^K�g�od�vi��	;���C?�`���2-w��W7�.�9b��4�x��io��շ<鈼����';���Mi��9�O�K�©y;.auwڽ]���(S��go��g�h��'��#��#~iGK�9����wT:Z
���5?�O=�$�����`�9��ݱ�晻#v,zFW�U��[K=���qӷ�F�M V��sH=�1R7�C�3�p�F�K�z�َ!�d��Xo~��-ѝ*zP�o�0�<g�;a�ck(s��f�I������5��}��m%1�QK��2!$��OT���t��4�P�?�6����fS�:P����X��ANtac��X�A㍳�T�o�'³�_�Pc�ݚ��hIm�E�;9�x�tb$=��oG���@>�Wez5ٺ�a-zMLn��8��~5����P*� S�{�k�]��F�ÜD�,�Ʉ	�֫�^h�U�����!:gp>K�ʕQ���U_���"����.��p�h��	\t4V�J|�|�Rh칕5cDl��*'�Lp�;�r���I��e�=���ʖ=����SN�k�x��1_��
�R)V,W�j�T������.l����e�-Vi�~��,ntԠm�(�e��չ�`��|�|�:%����Z����7�l�@ݚ�_��nr���������tw7ƒ(D�5��jn҂��u)4ѹ��(J��i=�h&[Bӣ���/�5u7�n�I�3@d/��A7�\I�tϗ��54��xS�`�#���^�^	�OӃ�o$|�������NZԂ���;GhA�#	u0�{��m�OM#؈>IA�L?_����7�+��.|��uѲ��O�zRW�Ȫ	Ww��v+�T�-> ����wQ���T���B�r�A�V,�-tGW���?@V�T�	��@)���z1����v`������d��t���5T��Xpל���4���`�3���P��*y���r��d���B߃N��}8�<-�j"�?�|RX��Ox�p���c秿f�ǭ��_������N�=�����S�Ni����^5E����܇�=iG��������2M`��9-U��� )�1����� �Hz�Ҙ)[�����U
�O?�]G�HX�MP���YA���h$�� �N�m�c5�NPG�e�_��kU~Ƚ�B�<�fn��j+#0��隁��4#���������2rMV�R,}N�#Ա�y�m�%K�m�N��I붛\4�ԓB�:B��Rt���=zy�s�r�N����2�j�pw
�_�ײ�fk�|��EAt�ʸ��kdW���=*gs�_��zӶF_I~*��Ze���{W��0\N�#˛�6���"�������3��ٶ}�F����.�٬a\Pwo!�OҾM|K��0V��8��ݤ���Kb���*_V���GR�,q/���e��ef7�sbdǪ *G�\O�qQ'���������[�vB�<3�A�ӂ�����*�I2aE\P.i�j�s-�/ۼzF%l<o;>��̻��?T�����u� R/�y�US�1�?���PiΌ�]bX+�ݳ��"$�"��| �S E8�v.Q�vҰI��,U�Ts�;Ϭ�l�0�k����s]�pdf���uT�c�c�v[��0AªY�N(~<�i�KWk�Z�n���I��7-�UՀSI�W6׼�@�,�o\D�@�Ɇ�f�E���1�	p�S]v��E;�g�Է�����]��y�i���*Y�Рl��>�@�=��k��;+c�țg�la�l�\|�Z�>�~�'ե��<9��*�%��܁�D+)υ|A�%�4�[
Mv�x��4�h�

5Ĝ���x�xx^�d�ﱳ�����f����:���7A͞�2Ư ���같��Bh�nT;� pR8���и�A����C�Ñ��Q�Gr|$��mq�������3�	.�O��%�f���!'Y��"(����r,�8.�X1?���E���-����H����R��{lz(�K�6
Mc/2�$B�J�
0|����ЎX�Ƣq��*��1�n����y&�X�q"m��ֹ4S��swuo�=�������˼���f\o������z��}�Pe����Û
�z��9��W!�L�J曚<�{�鯆?����c&�B���r��4��aO�k���(�m��Q�UZS'��84x�f%���t?�����z�����໫R���Y�Ң�lR�$W�ʆ�7������^��rt'�r~�l�}����h����v�D<�X�p$ۃ�G�.�B�؆~m:ZWɳ-��ށ|��*ywW
��d�E�`�] ��}=�J.m��lP"��<��I��l[��^���r�Hp�{���G�Q�����8�.(�O��q*p����`� +�ԭ݇R&�w��(��i}�N��kʖQYoɺE����U��&��*���\zj���_vuٗ�/:Y��g/�C�NJ�='84�`��P�n�?8V�Yuٸ��)g�A�ۚ�.D~��<L*g� ]􎯫~)�eZK���O��QK� {Cs���'���J���B#��Y]H�)Pۭ�q�ʑ�bINP���D�ZZqKŏW'�t���-q �nK���OW�o��B���F�F���M�Ƙ���Y�g_3j�����j��A]�.�E��|!�@me"�W�7�������܁<�χ�* 	��f�������2�n�*u/��h9���f�lw	�$c=�تcRh���O���d	�k�%��Xh�_��3K�<$�2Z�v�]���n<��~i �(����������3|���2!g{i����X�54z�P��;F�ɳ�J���ە�����)�������cUT���*C���<<�#�P_������,Ǵ,]�ڤ}�P,'ZR��6�3'��jY�+=�X��`�������Z,_'���g@���A7�N_~�Y���$7(�˹��Rml�ܯ~fĜ�d냏И����X�f�ʜ����
��:�;Q��vP-��[��1��.��B�9_��=Y���^P`
���?%-<
;�cܭн�ۧ{���'{���w2��9kA�/g:rw��� v6�,�t�������u'���t%�iz�<�D�:s,*��2�����c�k�ph�~�i�	�u�˿�Ga-�Sڊ���A�?��?'�2�>�a�3y��<�ɝI&��S\�U��E���Ӗޙ;j�9��,gu76ֿ��3T�y���AF>c�)L�臭��"
*?D�Χ�/
+�7Aʫ"VѦ[�}�<�����4��n;��j�N		_r�N�SCet��+&,�	m����ү���Eu��Isq�O��t趨��Nn��@��/���@]�K����H�����k�f�'�M�c�!n��4��]�J�v�Qr��W"WM�zmkn�pbAl�i+�r~��Β��*���T��fO�I4w*O̲aw��Ҩ����p�)����Z���x=������X����ҙ�g�ϴZ�]���6�*�+o�3�.n��F}!��+�<z�2�4=^N"靖\+g�a�v���	ѭ������w��]U�nn�d�|��ׯJ�nSޡ5�C&t���p��~�H#��Q!
@k݅=R�Ғ
�������k������.��s���&�����"=��.�m@lO��w���hQZ\�*�a�q0.���#.��;�[6�w�%��@٣��>-8sT�sk'^E�G��5m��I�1��=*��B`�L!�G���i���_W��h�)�Z�����T>/Q}� 9,�S��M�
9�T��t��Ab�gk��Mᯥ��CWg#!�t�Ϧ�)_����*�J�6���5��D^󇖴R�Ns���j|����l�9ۍ�tΟ����0.?+/��<b!��}Sd��"Ё�v�q��7��b#Rg�b*㕂JP/k���#B��<���Ⲳ�+4�W�X�ZK�uQ��������9���!�a���3�\�5�2&U9-���'0o�3�,�]I�Y�|��l��*|��-�l�YdkX�x���i�r�G�F<�i���})�Rtϼ'ѡs�m==Џ��\E�A_h=�A�E��t�Ji�mLO���1�'���F���V����𬰮O��{��3Ⱦ�:zFS%�����=�4��Bٝ����J�����p݅�G�򵎷�܂�?@\~Ai")gi䪘���n��i�F��%K�Z���tb\4��Q�xu�9râ#��",��T�q{�ً!�XE��]h\[x��� ԕ\�O5�~"=+�s`�R8n�Y�xz-���2O�h����1]��uA�-���Ȏ�����3����7���z��Mi�;�*���o-]��ˈ����[�����[�좼ݺ��~6#��\�um�WZ2sA� J�#���Dťg�*�Ɓ���W� ��L�Z7�it��t�N����c���rR�����Z'\��Ljk��k��?Kؘ�,r���T�U�ڻ��U]�֣����3�4�w��!���r��H�Wû s���B֝�Fk�q�9����ڻ��$�8N�Z�i��͝�nJ��y�H��6D:Xt��$���LG�h�m]�mI=(z�`M�,^�B)w�3�R�����0i� f��%�������v����=�����������}� m���Y��ŏ\�Gֆ�e�E�j*�4���I[e�����B�g�|�}���<�0\����ߥ��R�"���i�X;Y'���Q!V�tܼ�'Eq�ڸ�bx����t�;��v�?���H�4�������M�p �������ܕ*�V.�ʩ���J/z�י/1�S�������.��5�2��F19����<2�o]��*��S�ǆ`X�o=��Hd�܍ELV~b��7U5ͽM��9
!��Y�����VM����=ZR[�R�5��\_Q�Ύ�������"�����(I-�oE�G�.E���6��6�I��ȁ�Z��B�!S��)��n0!��=��#�5DL��>�o��%ĨϸG�h]�.L&(�Z⛕c_�UZw+�6d�DΝ5��@����G��đoj�@J�/Dm��+:���o1Z rE��LqZ��Y��G�[U� -Ab\�+�f�T�GK�����l�9b��
�%����4�n'6�*�%�Ax�Q�Q�4��N��w�q���V˾yf�Ynfg���+]��r��g�f�wۚ7��#X"%m2�jk���I�B�>ss[vr<gKO�.O���7	f���ToK[W���N	����&� ��sˌX��G\�T�m�ǵ 9 Oy��<�9a��$nS��Y&�>�X7};>�NȪx�����"��I`��%;m*1�-���D:M-{������Ъ�,����6Ǟ�NޟZ&5��1,�;n���/M?p��`NwqCQ�e�����R�ZFJ�8o�m�xYTϧ��3��4���S��1	���N���CC���=2	0 ��,K�
�6�9���O?R���z�x��E2���������PX� kY��w��RCxL[�P��ܥ������"e���ke11M�v���t���SP\pު�N��=��A�1�ʘ�jsd�^5�{�o;��9%g���^핯l�i�%�|�;8���]�d�h�_�N s�bC�Vn��(I���LbG#���{x=U?3"�t_iOm�ԧ��G(�y=�B�﵍R��v�u���	�&�R�^.FV����������ib�쯬����j�SS����q�c@�R�u�h��B�>Wj�"ҽ�>���9�X�|d����{J��] D6Z��Ƿشם�L�P���-~�	D���0B���3\xc���ɴd!�D�������Q��U�z !AB�� !AB���iԷ���T=W���� ����!B��k��;r�w
-��M�I��;>ߋ��Ye�,J���.�ݳs��܄��V�Z��G���'������C͂B!��E�ԪG�`���ιL�<�s� 'ՓI?v�&�b�"N&��Ѱr��(��%��^4W����*خ���`m3+��e�ë�8Mje�Ū�8�scl�Ӳ �ˌ:z�rȋ]l�}�@��('�<�5�H�;,���nl�D����XT��K�*؟�纳�Lc�`�l�l�\ _��m�e����9ѓ�o.��KްMeMs��,��t0���y�86���`�VLq�}��|_P״5�p���>$| �L��PK   {c�X�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   {c�X1���-  P     jsons/user_defined.json�\io��+l@=��з�do��-ER� ����&��hy��Y�O5I]�pFVd1�Dg�Uw�W]�`����M���8�1�4��0:�g�q5�/p�KW�K�o�����݇�:?{YM���]����+�5:[.n��ѧ������d'�x0��G.����k�P4�!��FªD�P�)�}�~6�Y�{�~>���c�tiK8�AEd�$�p,w�zʛ�gx�f<=��jt�[~��r:�y	��'�r1�}0������y5g���	\�J��+M`r�n���t"��\K"������R� ht��-a&&����BF��v��v����6Wnjve�*�|���a������fb�U���,aYV8_]T��+"J����Z��źI���nf�M�-�m�7_��t}3���e��	�O0#�͒�nϦG��ͽϙ]��qF��6�?/ǳL�<�yR���t��_,gq���`�l9^'Ӱ�π������W�5_�"��%X ��@�px'�2̙���N5����;Y�tm?��
����N~���+=���ä���\[:=�na��2]ss�R�'^jd3(&��� .�a�$I��Rţ�NG׈'Α!� 1}����L܌�a����DLa��%p�;
�N\bͭ�mj��'¯L��lYR�(_[h�7O�G�$%�Z�`r���=
�ǟ�v�!h� F�U�jś h[�����ZNC#�c(U*j�: �JR��@|8j4�w��%�F@ c��|�u��yi���J���7?�V��!Nޮ��v���S�uyWլx�����A�ŝ�?m���h"8�8��"�:	�q�+�3�НA���u�a!�� �E��f8�઩	_:���qj=r�HAj�H�J��§�4�;�4U2x��ʧ��3���g]r�.����;�7���������ίӣ�V7�iA䯴8�Gݲ�Gۈ�Np�r�Kdi�1ː"V
�<�^uN��p3��a��i"��!f��)����Ism��̓k�����c"�K�}Tڥof#%7�!A�%Q���l�b�AZ@|a�֢���N{��޺YY��y�.���}ܛ�Dge��=�?5G����`�d�\�g�J�~O�W�U`�+�����+1h#� �DB�0x'uB)�I������yC)X`HSH�8�5�%`哏ޤ���$-u����{��f}[{a�_��C���Vgnj�f�-v�rfW5DKȍ�N�C�R�h1�����An��(���*@/]Y�M	%$T!#5���!��j5�\�T���W�ɩ�Hd�a�c,A>��J�E0IJ=_��U�PA�M��(J��@�[<�V�O�*��#iU*��ɨ,�Nyd�qL��1Am�rZ���.���,N��Z�Sq;^|)���z5r��iKxw7�ǎ�*��˄d�0 1� ��w�D�Q�ո|�A=�/��4"��ư�sou-%*@1
���FA:��~|p |'���)���qw'�z�IK���o��(d���tmmD�G��>�SϚ�o��o�u&��u��B�k0�%�7vdm��_rG�ɠ@��1A �9Q���������bTP�3-:�M6�@�wI�������7D���x�u��C(����[�_��~-^�j	����! -�"������l�ʽ�@��l��筬xj�`�&㛣;�\�b���D�z������>��hR=��ޭ^�ƴ��ٍ�OEz�ʳ]�
��^�R5]\��9��a�#G��;+>��6g�l��I������<��
�\�9�(��n���=z�<�y���Aσ�=z�<�y���Aσ�=z�<�y���Aσ�=z�<�y��K�����1�8�nI�d��G@a�
)�VF}B�a�B z�򱫢%��G���@Z�D$X	�"��qB��qdx4�s#�!B��#��1*���V3\2��(���--t�{
��?k�h���[*ۧ����}G?���k .��?�<��) ���@8�<��g����s]N.�֣Ռ� ��V� �@� �u���jP5 �и; +���7l�z�z{y�h��,��E�E�M㢨Rq��1oY�����Y�$��%�@��J/;��HBl4yL�$�G�,�I��mM�H�A���Ni�)��er��-�/�$Ǆ\���C+�$��Y�2Qj��,FY)%�{:��~��%�{I5��Z�o����5�T/���h����p)�3ޫ3�@i�Uѧ;V�:z������{���-� S}ց6ϒ�#d-Hip�u�����$g��T����r�L��4���%�� �}�@��D��z��j���K�.��5��m{8ّ��:����G�ֈP5���~ �́�]:�.{��2I;�u�f�thY���dU���ꟸ`��W\�Lʮ m ;���a��<�c��3t��Wd�RM0� n6���
XB��t3���Qi�����6ݱ?S�K� ��N�f���3���P�u&Q@]�F�R(!�s�9^Ӻ�5�?'Ru��q��u+�~�T��Ӳ�uK�}"����5�K���C��:Ӈ}d/ں~��q�Ţ�v:�y|����D����Q�(�,Q!��R"&g��Z��|�t@�i0�1�;��2b9�ѱ��Ǔ�,wU)PCb���^���2w�1"���������u�Z��	e�	�����C�W�L�^�<g,t�r�~�W����S�-N�]��m�7�����Cq<��"Fq�!h���P�|\�bBB�-�����~��?PK
   {c�Xx��\�  oa                  cirkitFile.jsonPK
   {c�X��_�  >  /               images/17d126d1-8a97-48c5-9cdb-beb53ba7b71c.pngPK
   )_�X�C��z �� /             �8  images/182aae98-c01f-41d5-bd55-0eb3a1cf7144.pngPK
   {c�X��g  n  /             5� images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.pngPK
   {c�X����7  �  /             �� images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   {c�X����	  P  /             m� images/471995ad-a105-47c5-9945-45370623043a.pngPK
   {c�XhT���� ċ /             v� images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.pngPK
   (_�X��D>  ?>  /             I� images/61ab5d34-94e9-4496-9157-f8e280b3269a.pngPK
   *_�X� ��! �3 /             �� images/646dce44-14bb-4c05-881a-5e107587e346.pngPK
   {c�X�l��A Ԥ /             �� images/670050b8-4f2c-4603-900e-28b8075f4ca8.pngPK
   �m\XvO�XM�  Ի  /             K7 images/6bcbb164-c8eb-42ac-bbc5-5fd68c68ea6c.pngPK
   )_�XR�/�+ �/ /             �� images/74eaab8e-d748-4f44-9179-11cdc4bcdf9e.pngPK
   (_�X�����"  �"  /             �
 images/83968c91-e49e-422b-be2f-46fb404d4a04.pngPK
   '_�X��iP  K  /             ?
 images/8489a8f8-4880-44ba-919e-53c698ce78bf.pngPK
   {c�X�1.:�  )  /             �L
 images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK
   �m\X��>}��  .�  /             �k
 images/8ddf307d-15d9-469f-99e7-c830f4f75d99.pngPK
   {c�X�&�}[  y`  /             �[ images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   {c�X?S��� 2� /             �� images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   {c�X$�8�l  �  /             �� images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   '_�XF&�!    /             U� images/aa671e02-30c2-45f8-acb2-14f46084a715.pngPK
   '_�X����?  [G  /             �� images/c05be033-d934-4815-858b-3a150ff9d8b3.pngPK
   {c�X���لO  �� /             � images/cd9a76b9-8a14-4d7e-9261-140514b5ac3d.pngPK
   {c�X�GDU7� �� /             �[ images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK
   {c�X1���-  P               ? jsons/user_defined.jsonPK      �  jJ   